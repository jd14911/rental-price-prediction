��o       �builtins��getattr����keras.src.models.sequential��
Sequential����_unpickle_model���R��_io��BytesIO���)��B@� PK       ! +�M^?   ?      metadata.json{"keras_version": "3.6.0", "date_saved": "2025-01-06@14:01:17"}PK       ! t-xү  �     config.json{"module": "keras", "class_name": "Sequential", "config": {"name": "sequential_9", "trainable": true, "dtype": {"module": "keras", "class_name": "DTypePolicy", "config": {"name": "float32"}, "registered_name": null, "shared_object_id": 2309670233904}, "layers": [{"module": "keras.layers", "class_name": "InputLayer", "config": {"batch_shape": [null, 10], "dtype": "float32", "sparse": false, "name": "input_layer_9"}, "registered_name": null}, {"module": "keras.layers", "class_name": "Dense", "config": {"name": "dense_31", "trainable": true, "dtype": {"module": "keras", "class_name": "DTypePolicy", "config": {"name": "float32"}, "registered_name": null}, "units": 128, "activation": "relu", "use_bias": true, "kernel_initializer": {"module": "keras.initializers", "class_name": "GlorotUniform", "config": {"seed": null}, "registered_name": null}, "bias_initializer": {"module": "keras.initializers", "class_name": "Zeros", "config": {}, "registered_name": null}, "kernel_regularizer": {"module": "keras.regularizers", "class_name": "L2", "config": {"l2": 0.01}, "registered_name": null}, "bias_regularizer": null, "kernel_constraint": null, "bias_constraint": null}, "registered_name": null, "build_config": {"input_shape": [null, 10]}}, {"module": "keras.layers", "class_name": "Dropout", "config": {"name": "dropout_8", "trainable": true, "dtype": {"module": "keras", "class_name": "DTypePolicy", "config": {"name": "float32"}, "registered_name": null, "shared_object_id": 2309670233904}, "rate": 0.2, "seed": null, "noise_shape": null}, "registered_name": null}, {"module": "keras.layers", "class_name": "Dense", "config": {"name": "dense_32", "trainable": true, "dtype": {"module": "keras", "class_name": "DTypePolicy", "config": {"name": "float32"}, "registered_name": null, "shared_object_id": 2309670233904}, "units": 64, "activation": "relu", "use_bias": true, "kernel_initializer": {"module": "keras.initializers", "class_name": "GlorotUniform", "config": {"seed": null}, "registered_name": null}, "bias_initializer": {"module": "keras.initializers", "class_name": "Zeros", "config": {}, "registered_name": null}, "kernel_regularizer": {"module": "keras.regularizers", "class_name": "L2", "config": {"l2": 0.01}, "registered_name": null}, "bias_regularizer": null, "kernel_constraint": null, "bias_constraint": null}, "registered_name": null, "build_config": {"input_shape": [null, 128]}}, {"module": "keras.layers", "class_name": "Dropout", "config": {"name": "dropout_9", "trainable": true, "dtype": {"module": "keras", "class_name": "DTypePolicy", "config": {"name": "float32"}, "registered_name": null, "shared_object_id": 2309670233904}, "rate": 0.2, "seed": null, "noise_shape": null}, "registered_name": null}, {"module": "keras.layers", "class_name": "Dense", "config": {"name": "dense_33", "trainable": true, "dtype": {"module": "keras", "class_name": "DTypePolicy", "config": {"name": "float32"}, "registered_name": null, "shared_object_id": 2309670233904}, "units": 32, "activation": "relu", "use_bias": true, "kernel_initializer": {"module": "keras.initializers", "class_name": "GlorotUniform", "config": {"seed": null}, "registered_name": null}, "bias_initializer": {"module": "keras.initializers", "class_name": "Zeros", "config": {}, "registered_name": null}, "kernel_regularizer": {"module": "keras.regularizers", "class_name": "L2", "config": {"l2": 0.01}, "registered_name": null}, "bias_regularizer": null, "kernel_constraint": null, "bias_constraint": null}, "registered_name": null, "build_config": {"input_shape": [null, 64]}}, {"module": "keras.layers", "class_name": "Dense", "config": {"name": "dense_34", "trainable": true, "dtype": {"module": "keras", "class_name": "DTypePolicy", "config": {"name": "float32"}, "registered_name": null, "shared_object_id": 2309670233904}, "units": 1, "activation": "linear", "use_bias": true, "kernel_initializer": {"module": "keras.initializers", "class_name": "GlorotUniform", "config": {"seed": null}, "registered_name": null}, "bias_initializer": {"module": "keras.initializers", "class_name": "Zeros", "config": {}, "registered_name": null}, "kernel_regularizer": null, "bias_regularizer": null, "kernel_constraint": null, "bias_constraint": null}, "registered_name": null, "build_config": {"input_shape": [null, 32]}}], "build_input_shape": [null, 10]}, "registered_name": null, "build_config": {"input_shape": [null, 10]}, "compile_config": {"optimizer": {"module": "keras.optimizers", "class_name": "Adam", "config": {"name": "adam", "learning_rate": 0.0010000000474974513, "weight_decay": null, "clipnorm": null, "global_clipnorm": null, "clipvalue": null, "use_ema": false, "ema_momentum": 0.99, "ema_overwrite_frequency": null, "loss_scale_factor": null, "gradient_accumulation_steps": null, "beta_1": 0.9, "beta_2": 0.999, "epsilon": 1e-07, "amsgrad": false}, "registered_name": null}, "loss": "mean_absolute_error", "loss_weights": null, "metrics": null, "weighted_metrics": null, "run_eagerly": false, "steps_per_execution": 1, "jit_compile": false}}PK     (p&Z�n�� �    model.weights.h5�HDF

                    ���������     ��������        `              �       �                        �       �      TREE   ����������������        �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             HEAP    X       (       �              vars    layers  optimizer              0                                                         (      `       TREE    ����������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        HEAP    X              �                     P                                                                       SNOD         �             �      �             $            L     l                          H      h                                                                                                                                                                                                                    H      h       @         name                               �         GCOL                        sequential_9                  dense_31       	       dropout_8                     dense_32       	       dropout_9                     dense_33              dense_34              adam                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            �      �      TREE   ����������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                      HEAP    X       @       �              dense   dropout dense_1 dropout_1       dense_2 dense_3                                         p      �      TREE   ����������������        !                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             HEAP    X              �              vars           H                                                               SNOD         H             p      �             HC             pC      �E      0        �             (�      H�      8                   8     X             <             H<      h>              ��              �       �                                                                                                        X"      `       TREE   ����������������        �7                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             HEAP    X              �               0       1              @                                                       SNOD         P             x      �                                                                                                                                                                                                                                                                                                     x      �        @         name                               �                      (          
       �       
       �                                            �#                     x                                                                                                                             ��;]�=���> Z�>V�>�߂>:>��>��A<Z2�Y�>ܒ�;Xs> �[=�2d<��
>��=Tm>���>�A
>�xK>�r��9Ӎ>db�=��>����E=�_D>��f<p>���=�3�>*v�>X��=�(�=Pއ�C>[R4>�>.��>wI>o�9>4��=mR�>Y��>���=c��>�M��9>a!k="�T>�
?1&=��F>n��>�]@?�m�>�r2=�N�=T�>�З>F��=Yߊ>e�>w>-?PD�>=d�>���\�8>�&�>��%>p�e>�s>�>�(�<ݡ?	��=�?�[}>�}�>�e�=[Ȇ>"�>C�xk4?k�=៼>�y�<c$A��>i��>�>BV�+��>T>A�>�T��V�:� O�>�%e>W�j;mW>�~>҄H>kG�=�.�>���<Q��>䈂>��t=72>~"=�>��8>o(?r>r�=Js�>�=>���>p�>��8�{��>�$�=��=I>�>�>~�O?�$m?9��?G��?�^:?	�?.�?�@�?�^W?�>���-?�?ec?�Dd?�Sy?�PG?Q�3?���?�?r�e?)�7?Z�k?>�v?U�#?>N�=?gz?�f,?���?��K?kWp?йL?5�F?�{q?wn<��W�?]�K?v%?u^t?��x?�Ӏ?w6(?�b?��+?��?�&O?UyE?��?�&?eS@?�]?�I\?V�:?RG?4e�?V!)?n�b?��6?6:?Q*?<bE?��;?[>?��U?��p?9�W?m�}�m�R?�#z?�h?>m?�l�?�V?��"?�܏?�vO?�X�?�?�L ?���?0�@?�f?pk ��ݒ?fj?�:�?
F?{_?\�X?T��?e?����.0?��|?C�c?y��?�.���.?��?,�r?Bh?�,p?�j7?��3?�3i?8?��?*E?�?�>J?+�Z?�%t?��n?�:�?7eU?�C?l�,?M�<? �?�:?�x�?�k�?�'R?��T?UD?)L\?V�#?��=�}���=*=Z�_<۟�=
�+>g��>m���~����ۼ&R-�k%*>����kE>L�6��s>�*%>�M=z:>��:>�)�?0>:�u<	~=d�4�4=E;�=.܃>V��>�u9>,D�=8	��0>.���|]����>ojs>6����k=q��=M�=���=8�Q��솽��_=v��ូ�=הb=��i��=D��<#�F�b��,���Z>�;���n>Œ�=�BL>����͸=�u>��w�ngT=F>(��3>�jo>��0��=*j>�4;��->�S=��G�B�>��H>ecI>͚�>G�K��Ї1�P�t�>(��="�;=y�t>��B=nv==�˽6�_Q߼PV�=m	*�3#Q>%��u�|=>�3>$>��>�)�wh>�_>�����e�=��=�u���xD=H1D<
\ǽe��BH�<�����B4>�ӥ>狺=�ݹ=���=�L���a�=2U>�����E>��P>�,���+Y>�b*=([�=���n����=����%��K����p���7D�Y����;�4=ʵ>0/>�:.��3�ң��,����+>fa��9��=g�3:�� >V��F[����=ɷf>��^=��!;Y�ļ�5S>X� �;zI���Ǯ�܀*=�>ֽ=E�=.3��n8��սin>��>�Y>?>�~=M��s@�=Ԝ<#h =3	=�H>{AϾj��ɱ*>��^�,�<<���)��=�u4>K�)>�,b����<�{�<lцF�+��p$�ʱ<\�@�{��V��<��*�����}_>N|<C >�5� z������S��xȇ�z�'>[*����:�R��Е�=0^�����=�	��>���=�z� ����l��W >��M<Kف��=S#=2��==�<�0(�v�=���7��=n�\�%YS��f�=��K=w1>K���#c��.�<�]?=.���Wz>��ƽ�</�����޽��N=�O�o�u��'/��0���J�����4>�}��S��>>Sؽ�$�>L�v����N]U��k@L�a�7���Ȳ�:����z�2��v|>��?�.�<���<f1؇���<VK
�A��<pT���������v#>��M��Q��:�>J���\����%$�>�g�<}$��peE<�T1�s�5<��i��)=�F��+�EP>�g�<-u9�w�<:@��6�>%5�����Z����>V�B�8ƼVk⽖�~��y�=1{Խ^�=꽸<��>Cy=:(���8�����$�(�FD��>i����Jн� �>F;~��'�>���yӆ=x�E=���<�ۖ<ql醗��>�.�	��>��Լw�c�Eڍ�}�?f�4�l_�|+�z�߽�3<
s��vȈ�����Q�K�b� �d<U�<�����ݽn�����B�?<R��f=�t�����oA � 'H�)�=�L������ ���Ã�4�;�����x�*.�>$��`��R ��;��*=�AZ�ŝ�;�>��m>[c�=�7оLER>��1�����}��~�V���7ż�15>=1�=�6�6��+E�>�Y���V4>��5�'>̥��"&�<��!��t>�� >�Gy=����B�S=Yl��
��>`������\�p�e���r�=b���2�B
ѻ�L�;��h=����=�Z�=3w�=�]��oLѽ�d�;<�Y��F[>4�Ϻ��>>}/>Y�?��<��#> p�<�S����^=�К<M�->ڞ=4�>+��=#�4>&r"�� >��q�g��o�>:h4<X~�=I�=�J�>47>�+�>>��=r�=�Ĺ�����ն���p��} ?e�6�GG��2:��I���$ڕ>ޭ�=F,��Lf>"�>��<�)�����@>>�n :�e� N�<���=�C��9B�[6ý�C<��o>��0=��+>�R�=h�p=9,����=�v4>�������=��#=YY>>F�>ɃN>7���>�����r�e%y��e�=�Ry��Ӽ�����d#"��~|<̩���0>��佧�<����5O>t��Ė�=hlK=��^�WC�<���<v鼰j�=��7;ד���}��9|�YƩ���(=H0����=��=�}�=Ȭǻ��.>�@��_���w[>����-�@=~"O=Xk8>ꓠ;j)=�>:���~=c�g=RA>ۆ>+۾
>�v�=h�l���F<�VX�o<���<(��;*
�x��f�)=�>5�=���K�<��"��p�9�.���� ��="̯����=)#�=�C=�u��d�{=2��A4�=��<�t��M�"�&>�%H=舽���"
T=���������`ե��L�=P�f=. 	>��=�}6>�	
�gU¼r��� ��g꽜8 ̋,= v@=cO�=AؽUE5=$�=(�λ�.>�S>��=�E�=���7�>@�=ޓ��@�=!�˽��=���7>U��IV����<�v̽Ft�=:�A>}��=�b<���̬��w=��6=�8��.�o>���5���%>�L��I&)<l�^떵<'�ca�:��9��=����%>�8�=Y!��� =�ܓ;D��z�Y��ּU�ԽsP>�����=Dk�2Y��v#�<(d�����<��!���<��Qp=D�uB�=�N���)='I��Ac=�>�~�<A��h�߽7(�M>���Nʽ���(���P>��y��7>ӫ3>�)/=a�6�UmN�����<ü$��=���=�0�=~>�')��c����������Z7>��A=
o=��>�qn����=*L�<��i�k�v	��-�="�>w�!=>V<
�Ҿ���<#����=��=��彺���T���>M�������=ۤ˾�p���ۼJ��p�=(��=Ad�=��=�=sN�;ގ�=0�>:��<��=���=��Q��t�C>����=Z���b��=��=�c�N�f�2W<<[�R=�=����ŗ�˅(=ER=�E=�嫽�=>s�4>? �<�}���->�P�>�D=�t�>���=e����{Bc�->�\>k:>ȅq;d�V>��>t'�����=���=ة �⠢��*�<��b�G��ř߼���="^\>���>�e����z̹������>�E؇Ӌ�>����g4<���	d��T�=�H,>`D><s=>h�q>1Z��J"4<XK>�<f>�Vf=��r���=ؑ4>*�">�`���>4����"=7��=Dw|=���=R3>�V���-��6����<؅h#]�;���r'X>$긽���=6��<_>�'��I�=��|��IB=��v'�>=�ؼ�
�=N���X�L�3z�;)�>��F=�� > Nw����r��=�F�]���ig�<S��H�;?��	��u�=�K�J�>��=�����<��=*�=��@>
�	=�Yս�O>���=ɣ,>�u�=��^��s���=��x>�o��v+4>]�1>�O6>��0?xz��`_~>>E;���=�4>u��=�W�=D��=��='�#��/	>+�~=jAH>ۆ�=VT>>���KA����2ŰϽT�{�󆽧��=����(}�=^룻�φ�g�H�����8�c�=;�= F�U�d=��4����=/�#PB��F�<k�/� ��={�J��0;D��$ �=Y[��[I>0��=��c�$}	>>u������5�C�'<�*=�Η���9>��ؽY��;ޯ]<Ԃ�ưC>�4=]�Խ�9�dO�����I��`o<����m��u�=x>�69�?
=���F=���������=\/f��M>�� a=[t�=_��<M������=�%���><+��=F?��n��V<�|彴*�;)�'��|����=  e=hy�����_�B�g=C{Y��<>��Ԇ�J�=��>���"9�=R�=H��;�`����=qT!>L�	�9���{T���W���>5��=/��=ݹ3<؀���3 �N����d<>��.=���Y���/�=�S�����=�5<���=�V=SNOD         �"                                     9                                                                                                                                                                                                                                                                                                     �       �                                             :                     �                                                                                                                                             �B>�_>�5Ⱦ�;�>r>�>�Gc�>��1��Gg>F�P� GP>`z���D>?M?>�U>*DN>��>��K�Kw;�i>kzS>�:���gK><r]>�Ç>�0�|,�>n3/>�As>N���BE>�u>�p-�U��=H>�腼�s&�!�Q>�р>�M>�\`>��O>PX>Zc,>�V�>3e�>}��<<�>�K>U �>{�>���� 5>=�m>��M>w8)���\>pU>ĭ|>��>8<Q>X�>e>�ui>���5����H>a�m��d>�2B>�8>k�H>�]X>��v>bn>!���Gy>������j>�>$�D�b>-�=���b!�K!b>S~C��W>D�Z>��E>�1���c>���D�S>XC%=5�R�r�ҾC+�Pc>�JF>V�U>��'>�>�~^> �m>��U>ɛq>�N?�R�>�W>��a>��C>61#>s)2>�Ծ�Tm>�&i>UB�>�t�>��R>V<q>��ž�w$�m�x>d,y>`�<>:N>��>                  H<      h>      TREE   ����������������        �A                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             HEAP    X              �>              vars           H                                                                                 �B      `       TREE    ����������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        HEAP    X              HA                     P                                                                       SNOD         �>             ?      (A                                                                                                                                                                                                                                                                                                    ?      (A       @         name                            	   �                           pC      �E      TREE   ����������������        �H                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             HEAP    X              �E              vars           H                                                                                 J      `       TREE   ����������������        ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             HEAP    X              pH              0       1              @                                                       SNOD         F             0F      PH                                                                                                                                                                                                                                                                                                    0F      PH       @         name                               �                      (          �       @       �       @                                            �K       �              x                                                                                                                             �5�=��2>QZ ��L>9��=V�����2>�h��=�l>*3�h�=>�K�<}�%>O�8>�Ä>���=���=�E>��>�~>s��=G;>��#�b�">��[�K>z��=��q>H<^��o>��<U$�>�9�=ԐR>=49�;�=��U>e>�wl>��>m.�=��>��=�?�=��=C���,77&>v�!>˺�=��><=�=">,�0>d�=��<D;>9R�<[�#>=�d>)�t���[�T�s>1g@>�Z���>۸>g����u>^�,�<�c=�8'>��4�T�<L�9=g@��w8=	d>>�>�>>z��=\&=VR?>q#l>U�<>��F>!��P>;����+>N܀>h��=���f�?>��)=�k>X�>=��=p-���y>�w_<T��;@D8=� >�y1=��=将>�Q!>�4>H�7�چ8D�>�G>�M�=�D�= �>b>P�1>���=��=Q�>k@�<�>��>�I���4Y< q�>	f�>	n���>�Y�>�V'��>�5"�+�>��>���"��>Uy��	_��[�>��>�Ծ>sz�>���>Z��>�p�>%`�>ҫ�>���>T�7�>�>�a���>޼�>?��>R�^��[�>`N����>���>ي�>�d���>!c�>��>�Ģ>؃�>B�>q�>R��>�ҷ>��>�q����>�� ?^�>��>�=�>Ϡ�>���>8i�>Ɗ�D�>�?6��>D�>��F��>C�?ì�><̞�m[�>mu�>��	�Gj�>�m��{�>��>-c3����>�t����O~�>1i�>���>I�>�<�>c��>��>�X�>��>F��>96`�A�?ѰC���>m}�>�A�>�����>y/���b�>x��>X��>�"����>�� ?���>c��>�?���>��>�ĭ>�p�>4��>��;|ʰ�8��>��>6	�>s��>B��>���>���>+��>�����a�>$T�>B"�>{��>j��[��>�{g>��=nQL�'��<4 {>�b�7>�DQ�"�=B>��/��>y6[=�#�>��=��=ׇ�>�P>>S�><�>cP�=߹g>_�=�z>�凇S�={�3&s>�E.>��=M�>���9>X�=7��>`R�=X��=�g;>� m=��,=�r<��@>�zN>qV	>\�C>l?V>��>���y-v�=�=��>q��=,��=	�V>���=�,>��>��(<?��>��E>1��>��2=cI6��� >#�?�gw?א�\�h?t�a?dc�~�o?�P9�|j_?�P]?/��]?6�I���#�u]?�cn?��V?��s?�b�?�i? �t?�*M?�lV?�+n?�6�j�j?�L)���`?>'a?>yr?5��%X?^B�ڨx?�;n?N��?g/�W\?��o?	u?��^?\�o??Po?��?�vd?݅b?��[?�&�
��Uk?bGq?��`?Mh?�lb?1m?�h?�]?�����^?V{Y?p�j?��b?�܋�j?��=�5�=�I5>)�i>]s�k�= 3��v>� '>����?=I���+�:}F>�.[>o6>�՞>ƃ�=x@>�T�=u6>��>�>	���x�/>��&����=�8u>�c>5��"> e�m��<X}L>�Ӳ=�8�w>7>�;>��_>�x�,�,>�>u{�=�/�=�)�=4��=i�;�@y����=�sK>�=>r4S>ʂ�=�DP>�>�)n>���
�=l=�v6>��{>	�ćW��<1��?_r}?�{��Ib?��q?�jb"Vs?�����s?�t?f��M�l?���[�h?E�x?��h?e�l?�ۈ?��x?E�|?i7d?Ta?&uq?o�hMz?:�'T�t?1?`?^�q?�]Ӈ��c?a�佗�?�Pq?H�z?���;h?��?�ar?�{i?k3�?��q?�e�?�	�?O�l?NVs?xv?��b
�4r?�i?\?jwp?�3d?>Xt?%uh?��h?�ߔ��Gc?�t?CVy?ǚp?��.���}?h�>��1>~�s�T>从=9�x��1�=����u>��=�A(�p�;O=[�-��q>�(>�^/>��>���=�� >���=��Z>��>S�j>����>�haZ��=�5�=B�P>���"�=�����>$	=O�*>���>>�$>���=�f>M��=[Z�>.�0>���=�%n>�#=\�
I���>�_>�+>�X>�J>��;>=�)�7{�=	�<��P>RR|>�:'>gG>��>�oC�=�-��"$�����'�z���r�"�	^��8؇�����E�q�jY�]��j;�x&�Ԡ�#3�Ax����� 5ti�h����e�LǺ�!<z�ه�솆 ,����L���]<O5��*���!��a������(��зF�4��������2&�}���4�E��G`���-'�z����y\D�l[\�el��"��󳈇z7:K�-��
J�m.1��%1��ʗy��>R�.>�e�6�+>���=��]^>x���>8�U=��p�=+(?<0�@V�/>~i+>>H�=�4�=H�L>澣=2�~=O�I>�>o����O?>}݈���Y>�a>o�2>�S�Jm{>�Ļ݀�=�� >�k> ����3>A��=x>w"�=�>�N�=�]M>w]n>"++>@�0>8� ��`�	`>j�=�WX>t%�=�Œ>�W>�r�>�6�=b�C<b:~>�im>k�\>}�=� �V�=�#���ԏp��� ��X��Ǫ���臊(�,�x��T &�j�!�7( ,r"�O3��wk,c6ھ���`�2�T҇�\P� �+BЍA��]A�~�7�Qχ����DA�����T���B\Eg9� ���n,� e%���ڇJ�<]D��(6������쇸9n��(31�`3�R�3@2��_p܇��|�Z2�J�0�����4�dJ��߅�C������>��(>៲��e`>g�����5&7~>d��N�B	�=�T�=,G>�I#:����Z>E>k�=�R>`��=�Q>(�=�D�=v!�=P%z>r8���=8nq��;�AZ>vE�=w��0�s>Y�(=�	޻.��=�="���%j">�j�=T�C>��=��W>A>>F�=5w>�=
�>^����.!>�Aw>�p>��(>
��>���<�bH>p�<sݘ=��#>�;=8H�<�&�=�E<�\v�=Nw�=��1>}�%>�{W>���Sn=C��[>!��=�%��r>�|<Ȏχ�ʽ=��A>�v�>��=| >�	">�D�=��=EL�>���>��>@��"�	=b�>�E>��A1k�=��=ߏc=鐒=I�)>�F�,�>|����Y>��=���<�P-=� �=m�w>���>w9+>]�>��)��">gZ>�ь>?x�=OK6>�|�=�u7>&9�=]�)<
�=�}=�6�=�n�>�}���=n5>�#�=�eDX�=	'>�gh�E�*>0Y�]>xpJ>)_]]�=��=���i>��q>#��=�T>�8	>cB>Z�>>��=Ɲ�=[�&>�����E>�,U�3+8>z�.>b>����6>f�-=��=	�j>�+>̡����I>�\>�C>�>a��=��'>̓�=s�>�x>��6>Z���X>�r�=�.�=H4�=�G>��>8
�=ū>��=�D>3Jc>i�C> �=�M�̛C>*1C>[�=�φ��>�1Q>���t��:��)�(�<��=�v����=0b=ӹ����'>��=�zS>Je�=�w�=wT�
�=E�>��(> )B>ʶ<��=<��¤=�
.>��R>�t�Sr<E%=�4�=Vw?�=�w[��A>Vf�<�m+>i�><o�=��=r�]=��="_ >�pA=�
^��'��=�:>?=;�)>ʲ>1Z3>��>�o�=W��<�a�=���=nf"=��=�ll�M�I�$�w>�D=ץ���=<P>P9�nK>g
�r3>�
>�f��U_�<����<��>)��=Hu3>���<��(>؝�=q�>gm4>��f>���=涆�|>��ba$>>�x>Pf*>0����c>�5����<�[P>�B>���Y�=^N�=���=�!	=K��=l�">��=~�r>§l>�8>�B�u��9>��=�u>�rW>�9=>�t*>2ʋ>��S=X� ���O>��k>��>�L>]�!���=
͒?�H�?�q#��?���?_��0^�?�=�B�?��?^D�vU�?�WU���I�D�?��?��?���?�^�?��?[.�?)��?��y?cȋ?�V��0Q�?�?چ�q�?�m�?�ދ?K5�G��?�>����?�w�?���?�)8��O�?�Վ?�|�?�'?b�?�b�?1�?Z��?���?q��?h7�����F�?F@�?���?� �?��?W�?� �?���?Wۤ�
��?�·?ހ�?�8�?��5��?�z?��~?��h��md?��n?|l��{?�e3ww?<1s?�	�w_??g��v��"0m?+~?�e?��x?��?Bbm?��?zg?��d?�w}?�7'	Os?�i	�ku?:f?�~s? �E�%i?�/��	v?=d�?b��?��5_?Kd�?&2z?VZV?��?��u?fs�?��{?��h?��m?G��OV�i�r?��z?O�{?��_?k�e?f�l?[i?�nb?�-�F�i? �l?�}?���?�4���v?��>0�">�W%��F>+A>� ���;>���-�=��{>h��qD3>;v<����G>ҿ]>�Á>��>?ST>�_3>��v>dj+>�d>hL!>H�؆A3>����w|c>�>�}N>�M~��6{>�𪺮�+>7>�c>�&�����=�p>�>;[L>|�>�`I>~�6>��>��S>F�P>�MS���].>��v>*&:>T^>��Y>���>�>a>x��>0�j<Eχ> 3>�AN>dQ\>9ڝ��4�=���=��=�c�ڇ=[�3>�@�d�@>���9�>�
�=ɿ�¿W>��<t�1<�=��U>�@7>��>/�=��>`$�=*�=�'D=�i!>g7��W>H�DR>�o�=�g>�|��^��>:s<�ͽ=U;�<�/>Aņ�n��>M��=��>�G�=a�.>@�#>�D0>�J>��>V;M>-�C�"�@F>�U>�S�=112>���=�/O>\@>wu>��<n�D>�d�>�s>K��=��V>{Y�Ĭ�=p+�p��W��䫂ʶ4��^ͅ�CŇ��
�� �Ɔ�kD&1�����n��h�F�hBh%&b,�T� ���dk�)5�>�i\Hl ��˝"LD%n.h�b����>��&0tcQ�*����J*2������wL���?���
�0^��>M/(%U����)�p���
�B����&e��l@��������A:%(Q�D��Ў������q>>���=���b>f��=�o���>7&·2b�=og�>�9��q>�~(=���k=݈�=k��>�[>El>�>��>��>��=�t~>N���=���k�=��U>8��=g���+��>T�<|!1>԰�=_:|>��W�>�-�>�=�=�	l=(��=��=��">RS>�j�:��+=B����(��w>�	�>�7�=��s>�Ł>�> ��>��>l;=�5k>^�=J�9>IF;>�����=C��=iN'>pȅ��->4�>bɞ��kN>����5(>`��=)�����=�'�=l�<)>�y�=�2>z8>�*>o�>�2>�Q>�i>��>�і��C{>�킇^
A>��>�N�=d�m�.�?>	��<�O>��=�9}>�r<��>��>� �=_��=��7>q
9=��=�F>/aZ>8.>��Z.�\#>l��=�d>i�.>�8`>v>���=6>�=v�<>��> �>U�$>++��(�=?3>X�F>�*���=�c->ź�z�ڼC��<�
>3�!��S�=$l��ܪ�}>e�7>뜊>�WB>���=`}A>+>��+>L^z>Q)�= 0�S>���P�*>��=964>�|�g��=�<�;�B�>r�D>�y>�r	�3>/�P>{>2f>N�*>[�}>�=�H>�W>��=̺�ޤ��?�=�%>y�e>�B$>�(:>i�>h�=���>"��Uz>gH�=�S<)�=8쇨Ֆ=�k!���7��={�#��E�Tb��o�8��t��ܞ����)@���1�^m������� Mӄ��*�l��l�.[ـ��S�K/���$@��GІ̉�u�� �<�$;5�0�8ɇ����a��=�����,<�� 5�����+��:�J����~9�������8����X>�6�i����~���b8���:c;��o��՚��\q�\�v��be�QE����L�@R`�>_�=�ƪ��p>���>���� �B>�ޱ�SR>�\>�� �v�=:B8<!5@�HĖ=�n=>��W>Ŷc>B��=� >��=Z��=H�/>_W=Q_�
�=�Mw��f>r)>#E>'I��Jk>�t��3��=��>���=wV�0J>��=�=h�2>Mz�=׍�=��=��B>��_>ƃ=<���!�U�P>���<8�=�>ڬ >�m>�͋>��0>ۧ�<��'>M�]>�n>�/�=	��pQV=�2K>e<���-WB>j��;�Ў�9i>*�%�C8>��S>Ă���~>�o=��b>;z�>�N�>.�6>��=��>؀\>�0>�,>)��=Qp��	,�=!�9��u=���>G�	>S~+�=w=!`=�mn=�Y>!'>���gP�=��{=�h>W�	>��>?V�=�>�=���=c�B>J��<��$��I��ɇ=U˃>��{>��R>c4.>|�=�;Z>�~�=SQ=H>�ߑ>C[�>{n>``+�i�<
ċ>]?L>�=�� Q>�p>ߤT8I�=yb��>�.=�`�� �c>������$�V>91l>�3?>�|v>�	�=Y�F>3��= m%=	M>h
�>:̇�1�=h�Q�tD>�iX=�J>DP��&~>xXx�C>��=@/>�χ�}�=��=*C>Qr�=�f;>Q�<��=�s��n�<+c>�S�!�@�E>�=*>?� >םP>��;>C}U>u =���>���S?^>�%�=�d�=���>��1:>��t?o�b?�.�Ǣ`?��_?�����V?zb���_?"sL?�^��R?:x<����s�S?�4t?�zY?��`?��l?��a?k&s?Z/O???*j?���s�Y?V�?�u�X?�mO?:�d?���4U?6���h?�`?G_o?���V�A?۫e?�.b?ܢL?��d?�vU?Yq?�\?\iS?O?4���2U�_?&l?�MT?�H?��U?]a?!CM?pL?�Q�D?�`i?(�m?�X?��B�q?���=�>e�����==�+=B��_�<5'�=��N>(���Z>r'=n'g�+��=k�=�QW>��=�>���='x>:�R>~>3}1>���� �=��YQ�=��=�r>����� >3�+=�?>�:>���=8O�,�X<�]�<��=͗�=0�>6wQ>���=	��=kH>�=d�ɞӇ���=�b>Œ>>{�=�_>qŅ=��>0�s>)�=`>>�1(>&�>d����=�7>=qT>�7��O��=*��>��fP{>+�N,�>���=HS��>�;=慆�x̝>\�
>���>T��=��>K�`=��8><y�=㼂>�ݓ>���0">����1>>��<>B�w>���J�>~�=W��=, >DCd>�C1�5�>�$=�=>R5>�/�=��=�b6>)ȏ=;�#>��>��6����4>9�>Dw><�=>P��>�u�>?��>b�X>f�<��	>V�=��>-��>o?�@Ӄ>��>q��>5���'��>8��>��@��'�>�m�خ�>p��>ډ�s��>ө��wC����>3�>���>�Ͳ> �>e�>�n�>[��>2��>��>���N�>c-&��>�e�>���>&I�>4�y�e�>�Y�>Z�>��< ��>���>�>
N�>�>W��>���>{r�>:w�>x̜>�a(��*��>�S�>���>�h�>�H�>7#�>Hv�>���>E�h�W��>�G�>L��>��>��j�յ>��>/�>J&�L�=<�j>p���+�!>#z����?>��>���M�>B��!;>�P>vh0>�N�>��>�p>y��=@�>�N�=��>����5�>�p����=�o'>a�,>V��HL>cv���>��>��>f��K�= �&>�oE>>f >�3>�)>���=���=R��=J$�=\���FeA>�b>��M>@�>2�,>�#?>�kU=�`>ʘ�<ͥ>��$>��>=vx= � �}��<i?�=b�&>�<��-R�=�;>��c�0X>v�,) > >��|S`>q��<e��r�>�k>���>ͥC>���=ϙ=34�=�_>���=S��=�3j�> j�\�#>"C>��B>l����I>��3=��I>���<�N>�~���=Y�F�[w>nYB>��%>�%w>/>��>*F><�H>JP����4K�=D�=)#>I�>�->[��=@�=�\>L�<[2�=��>�� >��>�)��=�mj�,%��� !Ԇ��v���#��n
���υ��E�4���(�+�C���.��ͫV��x`���,�<ɇ�����Q.��<R��N3��k�24�|�>�������<i�ef��톇D��.�u/��&@�q�Lb��(0�m�5�$�p6�ݚ�&��|���<.���:����o-"=�N ����=	d��Q-����f<�I��Y'�z?��q?(M��0f?!�i?@^���n?�7>��fm?�Gl?,M�ng?X�G��@S�T?;�v?H�^?��m?r�?�Uf?��z?b?a?�[\?0�l?�`����d?e����o?�+`?��z?����h?�C�$Rv?,(l?e�?��6D&e?X�z?g?GRb?�Â?F#p?�G�?�2?�m?cgl?|g� |	��q?�At?�Of?�p`?Y0`?�n?��j?�_?69۽?M`?�h?or?�a?Z� ���|?���=.�U>��#Of�=�=!A<5b>iĖJۍ=rKi>\�v0>�r�;�� #��=6|�>�mV>�Sn><	>aw`>6?i=��m=�)=��.>�8Ǉ*:>�+���X>&Uz=�>s*��L�>2��<�ˏ=�>�LJ>���M>\�>�>>�ȣ=�d>ș=�� >���=T>��=>�[�`��W��=��@>�V>Q~�>�6m>���=-��>Rӻ=��=˄�=���=m��=��@=W*��">R�=�k#>��܇�>�v!>.ܪ�.�5=f:���k>�H>��чf8�=@j����\�p>��?>{ e>G#�=��=<r.>O>�=~1r>>f�8>��\DI>@���|�=���<+�D>�9���o>��(=�o>��^��=���A�>N��U�=|�*>�E>U�q>un�=W�7>�I�<g�>�S�3vY׷=e�
>Pń>�9�=(�> L>���QR>�k<��>^>r>�x>(�>i�և���=5qK>��>�Ũ4>��>��9�>o���cZ>C�w>2�����>>1{=��M�>z,>^�G>_�>�4>�z>�ր>I =}7�=M�b>�AǇ<C�=Km��$MK>{T{=�>W>���P(>W=^S>�ט>x�>rb(�a">H�<!�>z{>�B:>���=�$4>}/,>�D�>��>?P�=㧇Y�=��->#Ȕ>\b�>%�Q>F>�(>�%a>5�=qd�=�6>���=*F�>�m��<�=�P>��R�!	=\=:�ǅ(77>9����>{��=�Dt�<O���r��l8>&�>�֕>�C=��!>�>�/z=��g>"J�>/ϖ>����X�g>��h��_>5tr>��=���h� >{H;�fH>��>�2[>\N=��|>��>��"=�>Lf>�(�=��$>�/>�(>��G>��@�p��>W]>>X0f>��=6�;>�>2r>�4>����~�>N�%>S%>Q�=����o>	WI>��b>��4j>5�>����9>�u���=�[D>��r�l>�'�='����؈>w{�=�׌>�&8>�->s�f>��>��[>���=�>gHn���^>�~&��A>;�>�=��}�A>�O�=�>��2>% ->� ��(h>��}>�p�=�c�=��2>	+b=�};>qA�=��w>�_�>jX����h>�ei>w>Ecc>�)>�`�=��=֨�>��=ւ�>�r�>�W=>�y> a���;S>���=�p>�d�;�]�6>:�م�!�=v4�#?2>�7>HY��o0>t=�g3�0�:>mɋ=\�I>��X>�A�=f�=+,�=ʿ:pI;>W;>��x�<>�;�'?>��P>	�?>.ʆg�#>SWn<�.>r݊�y"�=�F&��<||T����=5��<��<{�o��n!�ۦ�==&>6Բ=�6Ň\���	�X>��=_˅>��b>��>@�>�>M��=((*<%=5>��=�>*>k�=E-J�=S>�s\>�|�=Cŀ=4���[>�O(�[��>\>�d'�Za�=W��=\؇GN>�a>�ب=�a>�V�=�>;�=ڰ�=�#�=��>"�wK>��L�0�.>� �=^>�yy�>4s�=�R4>5��>*��=F���?(>�yN>L��=��=�&.>{n�>-">��>N�>�y�=���9����=�P�=��W>Bփ>�Z>���=���=�>��f=`z=��H>��P>G�=NA8ȇ�=Ս�>�j->n�Y���>�VU>t�#E>�v�N>��=���{�=�����{��t9> ��=,��>X��=���=t�=7>�"u>�ȭ=�=U�ۇEe�=��j�/��=�N�>vHb>$� ���c>��<�>h�=��>P[�6�
>׫=���=�?o>���=*#B>^�>�jF=��`>D�	>�Kć�����V>��2>��f=�Yd>���>��>z�l>�>���<�3W>��=��>�>*�ɇ��2=���=�b->�XU>��>����� >a�Ǉ�>��m>��χ�r�=,��t����<=�ұ=C�>Z2~>|�>I�=� �=Kx&���=�N�=�
ּ=R���V)�=9ō>I�4>)����>R���h�;>V<��>���Щ�>�>�'h>"�'>��,>�Mr>���=Um[>�>�׵=�������>�&">�?">E�=)3�=yaf>�@>�A�>AE��r�=8�1>���=)o>A+h�ɐ=0�~>�rT>�U·p�>�t�>X-��X1>��o>*�>�u4��4>�_�=��/���>*��>I�>c�{>U�Q>bI�>qޥ>N�>̓�>�q�>n�u��d�># �ϟ�>Ŭ�>֚�>����d�>�P=5$�>���>k�x>����]>���>dX>��>�z�>��>X|>��7>�w>���>�C� z����>rk�>�~�>�D>G9�>�W�>�,q>X!e>�t�;��f>��B>3I>呢>�sξx>|�>��>�P���|8>h?�=-����/>/u���խ=0�2>݂ߙ�=\L�d�"���=�e>��2>�T@>�	>_�=s�>��->�Y�=JP�>�W��l>����e>F��=��W>����->��<l�">���={�W>��A��=\�%>�]>>�G>:��=E{>���=��=�;k=$�>���#�%�>�#>l>1�I>y�>�>*>/�{>�sp>��;�>�>�C>ٰ=�{��=ar>p*V>�/I[�>�9>f���J�0>G8�/>ʉ��M,� w�=�3+=D��,>��==��=e+T>���<%��=_e�=��)>�1�<ϙW>��l�>�}�D��=$qb;n\=�����d>��=@ =f�=P��=H#�{e>�1>�K�=�o[�I>>Dq�=eK[=�x6>>�>��U<�?��x�2w�c>�}�=p�=��=�W&>�*>��+==��=��O=��^>�ʈ>�:S=���=��ۅ����.=�^�='��Ԟ#=3�>��4���=K���>�se>��"�
M�=���<�Xf�|��=���=60U>�@^>�\>#�P>M�=(�+>.�F>u1_>�G��_>+�����N>xL>�>ߦ��`o>pb=�Q9>�n�<+>�^���/>9r�=�: >T5>��<A�J>�D�=�k�=�Q�<�fP>����Z��u��=�x>��x=�]>��>���>���<�p=�`;L~=��>z�	>�uw>B8y�>2u�=���>�%�~+Q=�O�=����~�>I�
M''>UcG>�.�?l>���6S��D>�'>^%�>@Ӆ>�>_��=�/>��=�X�>��v>�N���_>'dӇED>�=4V�=X�.>Z6>>[�;`�|>�&=K��>�}�u>��>�z�=�p>�>��-=z�>��{>�ӂ>��)>�^��D�Q�`{>�N�= ^D>և�>v�h>�9�=�%�=kxM>ۢ���xS>�#~>ɚK>+��>�����D�>xq�>�j�> "���>F�>���-�>.Z�J��>�ù>����>gh.�Y~$����>��>�{�>[��>��>+��>�O�>�h�>d�>B�>�	��,�>�ϡQ\�>�{�>͜>��Y�>{E��g��>Y��>�>�Y5�9�>��>��>�le>߱�>[�>z�>Z��>���>~�>��0�?J��	��>�S�>�1�>Q��>��>D�>��>H��>=Ȗ��>)4�>���>9��>���'�>"�=��f>+H4W��=���=ڸ���9>�#�C�=Vw�:����=!�T����o�=<��>m�>N�>\�>1�>6S>��=t��=0X=��
�G:>�:<�6�&>� D=��{>����>�~�=���=|�)>�yu9>Y$>�f;>��{>^��=��j>H�> &>n$3>F�A>��·LX���=��=ۑ>U�>�)>��p>x�C>F-5>;>���>F"8>��)>�3>gո�>���>פ}>��%�&�=���<�4J�Q�a=�A�Ml=�q><��_�'>}Ř:�,R�i�S>���=�%6=�S=>�G>5�$<�7D>~�=�L=|�=чa��<�uˇ��%>��m>�w>p��PJ�=��@�S��=��%>`xU>��B�kӨ=���=��=d0x=k�>�[e>��=y�%>�=y<;o>�ܪ��&!r>�Ay>|n�=c��=�e�=Ha�=0�=;��=�?�X>si>��<><_=����H>ۜ�=�̜>����c>Z�8>S����<7�#d�w=�c�=�H��7d;���f��-b>�`>��>D�>���=��=p1=�8�= :v>P(�;�Um�q�>�)9��>���>(��=��z���S>���;\��=��;>�Ѿ=Q�O��=X��;�B!=r�=�DD=Q}>��=c��=
s�<>����:���v>�H�=f�{>@č>v��>�=�I>�2�=�>ۼ�>+~�=���=��=�������=��?�`j?�D&��J?�}P?�Շ�z?^K�dYr?݅b?�bƆ+�d?�H�����5�Q?ʫt?eTj?i�d?�Yv?�?n?�p?�U?��c?� I?���o�d?��X��@_?6�B?6k?�,�U?��c��a`?��b?$�b?/�*���f?��x?5�\?�IS?��X?�}Z?��b?�u?�B?"�Z?����� �`?�[?D�N?)�d?�X\?�l?	 b?��L?$�)���P?�\?�Y_?.8n?ڷ��Q?M}�>�I>ӖR<9>�D>�0⇍K漰�+�>T�=��5>������c<!?�=��r���>*ѝ=D�>�>_>��A>*U>k��=!��=U��=.����x=R�4Mf>�b>�^C>�r��?�X<�*=#r*>j!�=�/>0�e��>�6�=&o,>&��jd>-�>	��=j��<J�;�\�=�����Bg=�f=^J�=�kS>��Z>0�>ِ>��>E< �3>ۜO>�:b>� >>V��m^>B�[>�3U>>�`ӱ[>g�O>�_�:
>�99�8%>A�=x�*�=ñ/<�=��2#>�o>��(>�o]>��%>"�>
>��V=�('>C}>5_k���>����>w[�>+�>��\�=0�F<3�V>�i>29>_�/[�i>n$�=~=�=q[B>�sR>��>m��=�@�=\�><�=��>�x*'�=>��s=R��=��;>�e�=��A>Gj�=hO7>z�:>>lO2>I�n=�/>��e7>�q�=�m=�����A=�OC>��ˇ�k>�Nˇ�>�D>�O@8��=�o��1���1>�k�=�2V>�h_>��=r=���=C5J>{�>��*>���]z=>H�%��=o�i>�f>"��{��=(#_��ف=@j[>�4>{��@c�<��9=N�>j=l>.��=�a>��>��=�c>�]>��ZH��HP>f>~Ԉ>���=�ӂ>ɼ\>uc�>[.B=�*�<��=Y��=�M}> �?>VC��no����=�]>�=��5^>`Ld>�|冽��=R��vB=q�@=�B����=����H�t��>�y�=A�b>fH	>�6>�\�=ܔ,>P��=�3�>weT>�����=?�K>P�>'=~>�Ŝp6>;8"��qX>��>>^�->�%2)�=�F>Vs >j�L>�]�=.|<>!ȋ=*=��>N2=H�m��mc>?�>j�>��>�qQ>��u>12q>Ƒ=�ȼ�\t>�։>zn�>'�Y>6�|;=�V>�*>eZN��y2>�H�<�8b*>�r�Z	J>
N�=�����4=鲝<nh:�|=�=��=y2A>��>�|�=�c>	n4=��F>e�A> �]=_8:��4T=&�ѧ�=h�=�4�=�W8��~�<��=�V>:��=���=Hr��tY>�}O=}�">��>1u<��q�<D��=m^=@��=0g�<
)����{�C�b1=�>��>�D�=bIM>\֒=�L>2��<�`�<���=���;��!<����+=��=tx>�,�3�>0l�=Ƈߨ�=�g=��I>��f>� � �=��� ��qm>�G/>�>t+�=p=5>O�p>�O�=�6>��=aO�>��B�ѱk> p���;C>9x�=��>uYL�h>C8�w��=4}>�o7>�ц�w>�}�=84�=^�\>�{H>u�7>�>���=0&O>���=w�)�甇257>
.>�>uy>\�T>���=��>�Վ>wL���	>hr>/E/>���>`�:dӏ>mv>���;��	,<|�u>�����=F��qUA>`��=� χ��>�9<��X��<�e*>���=~��=�/�=��d�=�4Q>�φ>
�=~,%�_~A>7�@�H>��>x
)>�և�\j>�=�p�=-/k>��8>L��o>�>�=�!�=�v�=~`>m/�=�=tɆ=:5���=Y�n�����=)��tF>q�7>$�=>��=��>��%>�]f:���;M+�>�=bD?>If=r��=�*0>�kx=(]2��<=|	>Tf��t,>L|*��b�=&�|>�s��4�=9�q=z���ݓ>z�>.�	>���=�~�=x'3>��>��>�9>t�/>�, �w��=�#�y>;m>>>��Շݯ>�6{=yA<��%>�O>����O)>�mc=A�=�y�=L>���=O��==��|�b=�[>P�n%I��Dz>�X=��@>a�>�Ek>:�6=8cT>j�>R��<خ4>��Y>ѯ=紷=�8�~�>�n.?��-?�5��(?�)?@Ԥ��6?��k���?��%?��8��?��R�є1d-?�o!?q�0?Q1?�2?��4?۹'?�e?!M'?�"?!��V�+?8p��.?�r?r�.?�Cj(?�o@��3? )?b-?�,����
?V�%?y]?Pe?!6?Y�&? �?%{$?N�?G�)? 'br!?F�?�
?�$?�Z*?��-?��?Ft*?�}���?b�!?�.?��<?�����,?o��>�k�>#���(>��>�����H>Kf2%�>qpz>+��X�>U�E=#�'��>��>x@Z>��->�TQ>��>��>��>A;>��">�$[�Hz�>�Eo��>j�$>,��>m#�>�I�<|x>���>G^�>��7��a�>i�>B��>���>���>j��>?>x`�>d�a>N>��6�@�±o>�RC>�TU>�qr>%��>�<{>y�>�>l�F�.r�>�
�=e��>�>p�/�>�pW=�	�=&����3>��=Fp,�����J�>�{>�{��,o>�|�=	[�=��.>�/>++>��=���<��>>Y=ݤ`>׷N<��!��=�C�<�>;�P>�T�=���r��=+��=��U>�;osc=&��� ($>Q�6>��>)'=�w>�P>�x�=�z=���=A�=�� ����t�=d�(>>�!e>�T>��v>���=�@
>�D*=��
=�b">مO>�^=	�&�5>N�^�9�S"��ߕEY ����r�bl��? �UH�^=�7�,�t{ƇB�B���
��X�]���* {$����E%5%'�f,<�O&:XXi�8���*�`4��) ��2h+��l��C����|��1� �'�[��P���L���W����$��O����+z��<�<��ґ^߿�ד��@mO0�=�6�\X�B�.����h�����O��p@�����>->ފ�B>\�l>��2>X�	��>�=-��=������=iA!�Q�����=�>s�2>7X�<��=/H�=��>�#B>Ÿ#>���=���U��=V���I�=�=Y>sZ��M<�&'��<>��=�u>��`��Y>�{�=�k>w@=�>>�w�=���=���h>�z>�0*�%3= �=SA(=0->t�>b�>���=;"�>/0c>	�V=���=!��>q�`=a�=&ʸ�xh��-#$>rV(>љJ��=���=�/e��>�7��{>��<��U ��=���<B_L�o f>1�=��>/$x>=�>$/	>�B�==T:�Ub=̾v>���;->�8�`�#>�]>�PA>��2�}��=hl<N�5�c�H=�.5>���> >+��<���=�>"�F>�b>�=��J>$q�=����2���]>��=BZ�=d�d=�T$>�^�>��a>�k�==���=�;g>�t|>� >DK�7AM>�r�=q>��u�<��=�Ȍ�2�=�	�vм<\Y>�&U� ��<,�=��FJ>K��=��X>�O�=���=�2>#�=$�=�'�='��=�M>���=����f;>�;�=�rM>[�և�^�=�>�<��!=��d�ET�=7�/M'f=G��=D��=fZq=�J >!�X>���=`�>�׉=R��=���Q<����=��s>��>#�>W(	>:�:>���=W,�=��<�o��*V>�f->��>�s:��;�><<&>��>��*[4�=Uу>�Ǉ�p�=\e	k�a;ǈ{>��z]�=^<Z߇�SI>��H>=�Z=���=�m>�<>?�#>�w>Zv]>\�>��·h3>�w��J�>>w�=�<>�&g����>qL<u�x>���=��/>?��\>�	Y>6�>���<U�R>n,�<²�=�Kj>'��=�;�=B���-�X/(>̛�=b/I>/� >~�^>a)F>��>v�>�Ė;��<>'��=KW>�N>㼙�S��=B�5=��>W���>>�sڇ���>����>n�+>ehP?k�=��b=�귇|>eQ�=J�>���=)NA>��P> �'>#�#>E>�>OCU>*�އ�>�qb�SV>Xt�=�am>�෇�do>Df�<a܀>.�+=}E>�����>_,�=���=X1>ڍ>�l�=ъ >S�>avd=�=>�ȉ������i>��>�gv>i`>��> pC>�8>?h|=XDJ=Qƿ=��>�z�>~ƒ>��R�=�)u>�->����akg>>ON>\ه���=����c >(�k>�x��#�=y���4?UX�(>n/�=�h>Zs<>�+>��\>�W>!�I>�5�=��D>��>x�.>���i]>HVi>�_>a�J5>�E��{!>}�>]�t>U��ee=�d�=�0o>Nn>�r4>��A>�G(>��=,��=��M>��;6�'�QA^>ǥ7>���=��X>��C>�z)>�:>�l">�~��c1>��>>(>:�A>����>��*>��>Q��?PK>rM�=G���}�>���J3>>r>0f�XP�<���ݓ��x>!>�>V��=TE.>��1>$��=n��=�[d>��=�@��ʺ;>f�<��A->��=���=�q�Q>���e�	>*D>��">P@��Gy>R�3>y�=A�=��=}>>1h�=>�,>�k�=I�&>|�3c�}>`ѽ=~�i>�W�=B;>h��=�;p>֍m>���ѡ=�M�=���<�20>TE(�3�o=t�Y?,�N?ZI�!H?�6R?��V�`�J?b�9��H?��B?��應�F?S�2��*�"}F?�)Y?�"L?�EQ?)dk?d�\?��X?:�A?�G?�D<?c�z�V?TކBWI?��G?��K?�e�EB?�d*�B�`?3�R?fc?�$ݱ:?s�U?B�A?�G?.�U?;eI?��`?Q?��>?�yR?�_Y�>[��<�P?�N?�RH?��@?+i??��U?�cD?��A?JA��zS?�ZX?|kU?"�S?0�)�X?W+>JpL=$��f�a>�k>T4��D>�K �!g>��6>�-·��>�6����]OH>y|�>p�>>b�>�>���=�g>@�>0�>�z>?�ʇaZ,>���4�O>V�@>��[><Ç��>�X�;��R>�_�=��^>�wX�>%y4>�O>�X�=��=�"x>�;>��M>�~�>m��=�S��=�����=Z^>8-1>�AU>��9>ӛR>.�Y>�À>m�<%b�=�7>+B>��>�����<�~�>��>�{�(�>��>����>Is�Af�>m��>k4����>�\���Ɔ���>��>C��>_�>^s�>��>ʶ�> �>:��>�[�>l����>ʮ"�t�>�;�>��>���>�>����I�>���>�5�>t&���>q!�>d��>;��>�Ư>��>%˹>u7�>L4�>[��>I���*�x�>'��>}��>��>k]�>OC�>ՙ�>�5�>�q��.�>���>6	�>�>�'���>u��>pE=;O��1�Q>�r>�)��=rņ��<D��=���Y�>��/=��CV�B>���=n��=�A=��x=�>VVf=0J[>O�=�T/>����3�=����r� <��x>r�>��Ѭl<���<�T4>�R�>z��=���^>��$>#�>�\=�0>7	>�΍=�0�=\�p>)�=�[%7��>1>���=��=cae>�^=���=p�=���=j�]�*�|>y�=),�=�:>ߡ܇�B*>FC2>��R>j5w�ҩI>7O�=9�,3�<�(t���=�I>'l�|�->sN�;1��`O	>Y�[=l��=��F>��=J��=�>�d=�1>a�>Ͻ�ǇT>'P��>�K�=tÒ=�t���	>�/L9ch>�\ >Aɩ=�����=�<=�Ș=�B\<:�&>	�f>Թ�=����(� >3�=�ׇ<���(i>?�.>�C?>4>�;>�r=��'=�n�=��W>�*$:B�'>j�h>�u�=a>���ـE>}<_?9�J?u6���$:?��`?�\�+�I?�����[?��=?��g�K5?*t����X�S?*�O?�W?9�5?ޛ_?��=?��G?F(:?��A?�T?�����RE?'� ��I?�:K?e�A?q�4��E?b�Ľp�T?�y;?B�Y?g�t�B?!�Z?�oY??�<?��W?�!6?G�V?��3?��6?�?Q?3B�����b�Y?[\I?�UM?�eG?�;O?o�Q?�@R?�|:?[aĽ9]>?j�I?C�W?�,3?�
��sM\?g��>HQ!>Ķ�]!>�w@>ڒ��/w�=��7�t>���=��lN>�&=�G��6R>�	>v&R>��H>���=�=(>5`>���;�>�\�<�&�ͥ_>�`ه��=��=T�>�.����=���� >T/>F�9>�%o��>̤�=���=�R�<�!>"2>i�>h��<?��=�%\>����	>=��=w5>|^K>=��=L�'>�p>y��=I*=8��<>ǘ4>ʁ�=��U��s>��7>��0><O��>t��>/*=��U>N��Wh>���=�	�
EC>l{�=��݇��b>C>�'U>q~>�C>�(�=��>��4>�E�>��\>��P\>(�C�6�:>���>��U>Q~���>�=%=ح�=��=�IF>����4>�>3�K>�$s>��>"l|>�xd>�f�=�4>��Z>��y�����>��j>销>C͎>:z�>I�>�2C>El%>_�<ֽ�=D�>X��>B\p>(d���>�M���a��54=g�7�Y�+��I���:/��P�%�2j�0e�(��Vq%�5��Q�>�t]+�d��~��@��I���'m98��)h#���l�@�,)���|�DA�{n.��s=�� ���*y��Ղ`5���(�(f� ˾� �t�|ew�$k��ч 2��@���G�yA1�b���@�M#���	F������CxĆ���l���6�ņ�B�m�h?�Fk?�5	��_Y?�I\?S��O�o?C'���f?p1`?�ْf�W?�u�|1���=e?��i?�)U?�nj?�0�?�D{?H�r?=;[?�zf?�m?�]�41q?�0��`?��c?�6l?�χWkh?�9K�6�z?{e?�}?�IUˢM?��w?KQj?N�Z?8�p?�zZ?G�|?Y?k�g?6�m?R�ʇ�̾_�g?�^l?�a?�]?0�f?3�i?=�j?Ҳh?%��H�[?�s?��r?�k?�)��d?�uO>���<@p�&|l>�Y�=e����1>d�P���>%�
> B%��b>���� ���S>�q>ޘ�>�=�	>�h>��=��M=��R>�<�=G{��6�H>i\��I>v>�>@�凎��=����ʠ=R>�b>��Ç���>İ.>�B8>��<>s�<>�?	>{|!>`�d>�/O>z�8>��.�~]N@�=���=<6b>!�I>7�Y>SD�=�~>W>��<�P=M>r�x>��a>�W�=>���V=�}�?B=x?��9�h?P�l?��τ�s?����t?��p?g��֭i?Z(���-��b?�n?vze?CMq?���?A�v?��}?21b?h�U?6�x?�6;.q?�u�P�b?ؙj?�o?���b�i?�����?I-z?���?4�U?�R�?�,�?�b?��{?Bzt?B$�?��p?#�c?��n?�]���h��2�u? Jz?�uh?��i?��f?��l?qw?�l?5\ýP�j?1i?|�u?2�y?0i�?T�_<1��=ͥ���L>�,g>�k���>/~t�=���=�H�#���=L����>��Z>^.>�<�U> P=#T=&>�z[>��B>J#%�=���>]�=N`|=� ���<�ȱ<��>��$>G��=#I@�j�P>��;>J��=���=�J>�V�>p�X=�4>��6>�N�=���$&��C�=�J=5��;n��=��=_�&>�>S(W>ޮ�<K&>8�I=�,>9qh=�U���TF���>��==P��P�@>��/>&橇�>f[/�UP;<"��==��a>f��<�j����:<�]>�1�=(`t>K�>�(>�1�=�g�=��G><�*=�几{L=�T:H�=��(>d��=vl�T�n>R(=$|8>�'>[��=v�)���<��B>?�>ي#>[�d>&�`>$�=��;�`>}d�=4Tw�sa��>�(>x�>�3|=C�=��G>��L>���=��3=(q>+"W>��b>h��=��wDo>�9>>W��=�	��C�I>�}P>&>��=Ⱦ݆Ѐc>K>F���&ň=��<Ͱ����=g��=��G>�7>`�=  W=�>u#>��=dډ<�ɘ� �>��as�=H�G>9�k>>qه��>�-���pi> V^=�.�=�f=�~�>��=�|>Ғ�=�>m=��Z>���=�8�=�,=���=�e'J�-+�N>�e�=�p�=~>z��=h>�GA>
� >jL�=A���/>��>�ɒ< �.+�>��]?f�_?�N?��Y?�����]?~2���R?~d^?`r�'�M?�H5��畇�S?�=`?�O?>>U?��u?��Z?�f?k�F?A5B?�Z\?n�;y�`?����O?�pO?�:^?r���̲S?\����X?�[?c�s?�z��pE?��e?��W?�HN?;g?�?N?jm?c7P?��H?�{W?����!K@�ua?�}_?;�O?��J?FW?��T?�P^?��G?R�ν$�a?YY?��[?3fa?��i(�i?�/>�=&|�H=a��;|Y�Yc>@��6N�=��=�Q@I��=�In=D��E�=��$=z�>)�[=t�=z�=�=�e1>כ>��<P=���h2=:��n�>Tc>�� >`a	>x߶<�}m��/>Ҩ�=p� u�=2(>x$%>�>W=���='Z`=��-<��=3Oa>��#>eJ���5��C¯=:5<$�=B�5>-�A>��A>sS?>8@�=��<%�=ÀB>�$q>?�4>c��(LF>Zu���������@`Їʬ:�R�ø�� ���$�t�����i��L�@����x��H���Щ��!���BL��t�ѵ��Bd��&�~�Z�����D���j��8��
�V� � �&����R��>����zE_�ڝVd2������;��{���&� 8R}��z��)�ȉ��.e�X�҇*F���xAfH)��:5����ذ<�loz��l��J(���>>��h=N`tY+>���=GWp���=��e��=��<#���s�=M�;VO3��=;6�>�b>��9>��!>^��=�Q6>�?>�+>h1 >Ň��	>Qׇ�\M>c�=�V�>�)�(�>��ܻ��=-\G>�]�=����p>_^4>r&>a��=�^>nm>N��=�1#>���=]�4=��8�m�4{>ӻ9>���=�� >�0>�
>q�2>L��=̽��zR>ʄ�>G�E>蹩=�:����=Cj�>Y�=>�RhVOz>��b>>+��1k>��B��>3d�>������p>�g�=,ׇ.~>}�/>Ч`>�>9\>��x>�H]>��;>)vB>*	>����G/>VbM�H> 4^>ia_>n�����x>���=*@�>���=�V>����n�>OJ�>�Hr>�m�=M!7>`��>Ii.>��>U8>��=xY)�;�:�K��=ηj>O>��>@ڃ>��K>23>wv\>|��=�� >�v>k��>g�9>@o��g=|��>�<�>6�)��mG>u�>��ꇦ0�>A�&<�g>���>p]�f�>2�<�K�i�>$��>Ox>ތ�>%�>���>���>	z�>1��>��i>V�2���>�\C�l�>0c�>�g�>�V_���>��;���>D4z>��>�>�*Ŕ>��>&��>ƭ�>�1�>��>G�>UtX>��>��>�����5��� �>Z��>�>Ds�>K֙>IzK>A��>�}>@ί;~ʩ>I��>e��>n׵>�IɆ��Z>��^?�kZ?@ԙ�|3?��=?��
��JX?]� �JS?�m\?�?����@?=x�C!��;?��M?&Y?J�5?��l?~�N?J�Z?Y�/?�(4?L�U?Pq��N?��ri�Y?�GL?LM\?356��@?3hc���g?4J?�Z?<�ZI�=?��\?�]f?��C?v�_?�:k?�T?�eB?��U?��S?D�@�{X0��'M?�Y?�N?@.X?B�D?��E?&�??CX?n�+���c?j?Z?�XM?�]F?�(؇��\?s,���͇�^`f�ʆI��7����=����� ��,>�{A������Y�����v¡?���v!��F���f�$��=F"��^7
�S�%�MZ�\��\�� ׅJ�e�%mD@�����@V>�����%��S���,{��u������v'&�����*:�����ˇ����&ć �J_�`�����E�0�.P�_�+�N?�H-;'1	�~�\���+>N���%;>se�=���$==���H�U>&��<I`ÇY��=��=t�X�9�>R
.>�F>��Ѽt}G��`=�P�=�?	>�f>o>�2�ud>��wy�=��y>� > 'W�Z�h=\۸<	�W>��[>��;˟Շ;s>�=$>��>Oj>\��=G(q>��Q;��<�弜-*<�\�I�(�0h�=�u�c�9>�\>�4C>&��<�ah<y�I>:�<^����=ql�=��>Q���k>J�˻�R$>��;Gp2>L�U>��d�>b�ml'>I��=H�0��=6�<����>�V�=��;8S=>Pj9=�n�=�R�=6�<��=b����`��=�-���=�Ul>U�q<���3M(>m��<�Ҽ�G�=!�=>��#��-p>-T�=��?�=��=���=J�=`B7= �<���=�c��q{>2�>�=��=��&>_�=D�2��0�=xU�<�m/>Uq>�SY>~>p>���8:=7�>�=��6\�=|������У>�X���	=�B�<�>�'=�X���>8.1>��=<�>?8>���<�"�=��=���<�E�>�$/?>Y>��=����=;�e>�7>���*>��`<��>@o�=?3�>Uz�>�DE���=��>fG�=y�~>�9K=��<̑=�7�==��s&�jQ=�$^>��~=�>\K>z��=(�u>BL>�N�<}�=>	>h�>�C>p��Ya>P�=���=pq��X;o>)X=�aǆ��>d��l>���=F����=;Aa<���N��=2�u>�*}>��a>z�>�!�=H�>(z<9L>��<>s��7@>�L���0>�tK>g�~>��i��^ >j��<��[=oiJ>_A>L���=g��<&�=�(8=�>	> �=e�>�Q>rd>(�/> ]�v@ׇ�>�a>[e>K��=�=��><�$>�>Үk<wgK>G]�=D�Q>�=N>�^�*��="
�=�1�>po�N�=�{>���B|��b�����8>�τ>��ܒ�=��2=��=<��=U�/>	��>��>��P>��=F�>-^�=_ɤ=�=���=�3��G�@>��4>�'�=�r�'Kn>t+=�>��h> ��=haN��>~u�=6>��=�B�=q�=ȓ>�ڇ>�0>�b=T��x<��~>��7>f>��>��.=<�2>ʉ�=i�d>{}�<���>�=���>�w=��͆�:�W�>B�>>)�)���A>��=��@�ew�=�"��#��=3_U>TR�i�=<��B�,�x_=m��<>�T>m<$;a��=cA>�"R>��>l�V>�t>��(���->��9�t�>�$>!V�={�)�D{>�x��Z`=�	s:KL8>L�>��>�FE>�!>�4K>ޡ.>��;>eY�=��C>��>]��;�:��ˤ���V>S"y>u�<>��J>�I>�W�=֓D>�=7"��:�=#�o>��k>r�:�`	�_�=�>�5r>񑍇�(c=���<uml�>�Vǆ4:=�h��z��$=	�;w6����=�%>��F>�i3>��u=}�=�qd=%F>pm�;~l>����@1=?���p�T>�;v<g�}>���k>���ʍ�>e�Y>�9>��X>:�;=�w�=8�!>�ͮ=fQ6>F��=��=i�=�9�=�6Ї�}1�a	>���<�>���=�Z=�->��3>N�=%$���#>�r>`kw>�z,><�>���=�^�=��_>4U��>�����>�g쇎	 >J�wu��=�=��^�
>W=D,���e�=�+=#�>)@�=�>�=�l8>¹�=�w8>:���:�~g=���A��=��,>��u>�W���b>@П<H�J>�>�7>�y����m>�?�;�I>:<>�j�=ߚ>���=鑌=�R�=��p>Bч�E��X�> �=�.>��K>���=8��=��#>F�m>��A<z7>��t>y>#S�<~< ��>9W">-�E>��l4�=��L>�1�Q@>�S �<�>Ѐ�=ܿ��rb�=�pҼ�����=ǘ�=AaR>�:>�/">�E���/>� b>,�d>	���|m�n��=�##I_%>A+�=Ā>y�">&�=@c�99H">�{$�W�>*w��� >�+>�pP=��B>�?>�E�=L��=��#>��=��O>�z��%iA�\_�>J�v>jC1>�ۅ>��k>%>��I>�-~>�$����=%�B>�Z�=���=to��n=�?(�?3�r�}�l?Z*q?3��De?P�9���o?C*u?�%e�(`?r�R�5+�m�l?�Ut?��n?$Lm?.V�?c�v?��w?�{\?y�a?�sm?�L��6v?�r���}m?K�j?'��?h+5���]?�����r?�Dw?���?����^?qZx?ݹr?�a?�Lx?��k?��?�{?��e?�y?w]:.��uk}?�|?��o?K:b?Y�o?��s?��r?�}Y?M�ݽl?`y?nxy?��u?������?R4K>0�_=�1��+�>އ;>/��ʹl=��@7Y>���=���� �=��?;�ⳇ;�!>��V= �=t�`=���=,Q>&^+>��=H�t>�	>���T|>D�u�h�=j�>h�&>���<�>i�=3=GL>���= �^�Z>��=�->x�Q>�
>}>`�=�I=�(l>G>0��6XC�=jaJ>��k>El;=�j>�k>]�>��=]�X�Q�/�D5>�.>��>xJ[���=�yo>��}>�v�	>�i�>N@�/��>���S�]>�k�>D@��(%>�R�=�ևw�=m=>Yp>�>Q>_�=�:<>ĒE>��=u�5>\��Z|�>���6>���>�l!>��̇Ǳ`>2�=��y>��v>Jm>nJ,g>�>f�!>	x#>�-�>*W�=��>���=��>��">�/�6�׎�>,^p>��[>�5>ҍ>�Ђ=��D>��\>L��<N�_>|��>��g>X&�>r%���|0>���>D>W�0���=
�='����> �5F�<5u�=��5�D-P>�D<B󇷷�=���=/>��>>�7>z��<�Y�=���=�:7=�h/>��Ї�#�<��i��=��2>	j>��D5?>�,�<-�4>�h�=z�=��]�=�2>��=�/>��:>85�=`>ҏ>>��>ĈS<�c-� �Kf>�_(>6��>06|=�6&>�m�=��a>Y#>��7;. >Jf[>8�,>��=��2�=8K>^��=��t���>(ߊ=����;ü:̶��J�=�&v>��)�c>H@=��=��\V>�䄻�>��<���=��9Ҥ=#�0=�V�=���>;��G	>6��>�C=��>$����=�B=Y>p�8�� >�m5���.<��e=�ͣ=�#<>Qv>��=���=I�J>��=� F>���B���=Pf�=��6>��'>7�>Qo> �;;ƴ=�>�8��>W�<>m�=�>+>+��{�<��>��i>�"��F=���>�ZL���=Pf����=��>��+�.u>��=�s��J8>ا�=��f>D�]>�uI>�>�W#>��w=�|t>��:>hX�.�>=���H�>5�>��c>����=>(CS=�Aw>�ҙ=�	�=���Q~=�0>v�>�h�<q�Z>�x->R�>u=�)>m�X>t���?��>ⱀ>�!�=<1$>UH7>	\�=��=PSy>��=2h6>=�>��>P�J>�i��Ch=�:�=PJ�>F9����=>�+>���e�=F��2> 6�>������M>�I�<�	oR=j�<>��%>�YM>R��=��W>Wt>�jV>_�=*l�=e
:�$�=T���t�=:��=kG@>Q"S�S�T>�����P>��=ت
>H��x(=0l�=�!>9	U>�6\>%`�="�5>3�=�fI>\��=ށ2��o���c>�'�=�ä>���= ��=�;>F�>f#>��;V�Y>�s1>CO>��=to���Q>T�?h�?�g��Z�>Ԥ?~u1��c�>4PJ���?�>�Q�d��>�+;�ӝR���>��>��?��?��>��?��?��>�y�>� �>8 #���>Ib�y�?�y�>�l?� ���?/��{\?Q��>�n?�����>˺�>�2?�I�>Hb�>a��>���>�A�>\��>�^�>}6� �F��>���>�h?c?@O�>t�
?�?n@?��a��Y?~?��?��>�v��?t�T>z/K>>��<�)k>mC��i=e�E�S=QLj>a����)>��<�~�ld>T�	>�`h>\�=ˮu=��>�o�=A��<��>10">�����=����">t�=C�>�Yˇ/T>�yS;:��=w8�=K��=QK����]>����خD>�->�=�1>>&�=iڼFJR>=�'=l�.��7����=
 �=�T�>�z>G�=?�->���=�i7>o�=J'��ec�=*&x>�"<�2��iZ>�g�>��>��6��j�=r��=LV �i�<�k�I�>/E�=�ކ�H%>ƭ�;����L�>�ݑ>�>��7>�">3�(=�)>iƖ=cWv>̔=b���
>�%7�e>-u>��=¾އ��>�/v<�,�<<1�>��>����� o>�d>-~>��d>��N>��0=��>��T>D>z>�t�=�Ё�?�>���=���=���=��o>�Wy>�ؿ=<w�=s��<�}>���>;��=l�P>�7և�%>��=G�>9�"l'�=錉>���['>I0�����>ъ9>n���Rk��I8��^%#>�>��\>�55>_�,>��}=��3>�u><>F�>����6j>s�i�`�>��d=by>�+��%K�>�-�bay>l>�t>�@h�>��g>��{=K4>��4>�7>�>Iw�>�՚=��2>�E�^�-k>H5�=�>V�>��	>,?�=x	>�>���<u�/>��>�j�=��g>i���tr>��=�N>�b܆$#>�\l>�+�'�=�G2�K�=MNo>���N>��|=Y����`><w�=�ε=�J>x>��=�p3>u~)>a~>��N>�b�v�d=��w��=>O�M>�o>j�ˇ2�>+��<L�=��F>�)>ݻ�g�!>��>�-�=d>���=��>�t>�%�=�O�=��=��a׽;�r�U>s83>]�}>�d�>s�>�]t>�<�=��e>��c<��.>��=K�*>�@>)!����>a�,>�yM=.��!�=�,�=�X�b5�=ד�OS�=���<�����k=��E=�Q�E�1=��6>)�_>w-�=g==��=Z>TE�;K��=o�:�۽��o�=����=��S>���=L��&L>�%!=�f>:;>z�>,�Kr>�z=!��<%^>��>=�z�=ig =!X>{]>Z�=&_�&�Qت=��j>U!>�+C>A�~>�"=�c��cx>Y��<�>;��=j@�=�k>G^H2=Fp>
�'>Dv��	>`X;>�o�c>�����>ů+>xY4��#>;��; .��Ka`>$�,>Q�@>	k�=�.>i1y=�>�=�ki>5�<��c>pc��/�=�n���=H">Y�v>����NS>n�=��<���<���=�PG7 C>n��<>�>>N|&=~�$>�9K>�=5p>p��=���=Ou�
�K>oA>ۄy>@̐>��*>�6.>�>��7>Q%���+�>�i�=2>
�>��!,=��c?"�P?�il�ZLE?vD?�r����]?wvï\?�:\?�I���F?�K���·�S?��`?[�`?*�e?��?�5`?��]?�YA?�M?�%M?JU܇Z�\?�����i_?�]Z?��_?k���ט\?�vB���S?��<?0i?��%�trC?`[?�`?�!U?Ev?3�f?:f?;M?�g?o�l?�C��VV�U?h�Q?��\?��h?�ZW?([?vBd?ccZ?��-���]?�`b?֭e?�{D?�O�R<Z?��L?!C?���6K?�(I?���YJ?d~܆��N?qH?��5�8?;����߆�K?��B?��F?��M?� [?&�R?Z�K?	<?N�<?�8J?m�$�vU?	��(�K?R�F?�>Q?�2�K�O?)� ���J?��M?~_?nw��-D?h_^?y�Z?}w??,�L?ίE?>�]?��A?U}E?Q"Y?o�������K?�T?f�F?}K?��B?ĭ\?�F?��=?���HA?T�L?��V?�C?细��P\?rD�>���>�4G���=��3>��>�<c�@�>PdS=����^7=��;�67 >�~>ش>:9�=�c�=���=���=�A�9ѳY>�tA>��;n�<�� ���>ʆ>��=[ �����==�;��W>���=��>ĉ���>�=�w>#f>�HI>b�}=��$>�*>�Ԇ>Y��=rJ��Qi���=��]=#E�=u��>�	>���=R�>�G>s�f�nƊ=��=�>Y�,>���NC&>�\�>'�>�`�[>';>������<3��4>w��=�ֈ�y��;�J[!>V�#>X8>+�B>~->hBc>��>�ъ=��g>��,>��X�6�<����� >��=O�i>F���K�> g��L��=��=�2>e]�u��=���>�� >�`L>���=�ӛ>~�>E�=��>�o>t(Ȇ� ��>o�_=R�\>:��==)>�n�=��m>�X�=�����7�=���=�a4>|>���3�f>�4>��0>�! �Z�;��S>��h�%>�0�T�,>�H�=��i��;>S=�9���!R>O��<)O>�?i>��=��=7x>__
>fF>��<۴��l8>H�j{n	>��N>��$>t���[Vx>�\�<��=�w�<y�=�\���GX=�_�=<r�=_<>Y��=���=�0�=�H>�_)>&U�=�9�?��Y>��V>:�#>�6�=q�`>#F>��}>R�>;��<\�8>�J�=6��=��Z<����=jϣ<�H�=�r����=o,F>�_Ƈ�_>� 0�?d�<~��=���)>|�<}Э��T>�<>�u#>U��<�%>�<��/>}�=�%�:�>G��oB=�.��f�=>��=�"��j>�Κ=�76>�[t>�
�=��3><S<=��o<!��={<�gW>c�=y�=P��=�6<7(.����&�=�Ky>�T>qz|>3;=;�>��c���5>���<�/M=���=aX�= B;=�4���Y>���=�n>�B�?�=�]I>�|���>��@",�=�1�=,/;���;׍=�'�C�>Ok�>�%y>��3>�DN>�j>�/>ѽ�=nS>�W>��	C`>�����>�pc>�B[>�ԇ�\�=��<�:>nZ@>!�>F�ۆ�[2>�w�<��!>7x:>�UB=x�E>r�=s`g=<x�=��9>�2	,T1�2>v*>��>�2�>�i>&�>�S�>�B>��<�#�=���=}�A>aM�=��	�k�=SNOD         pJ                                     ��                                                                                                                                                                                                                                                                                                     @       @                                            ��                     �                                                                                                                                             �G?��)?f��Pa?��"?bܺ�l�?H����?�; ?�����p"?�K���Ӽ}�"?�?��4?d�?Y�(?a�?��"?��?E�&?�p ?o4'���$?\��+�?��&?�3?�!��/&?`<���?1�?�M ?!�(���*?�?��?z"?��(?��"?W!?��?_�?�$?���B����!?��?�n-?`h-?&�0?�4?�?�8+?@�4�GI*?�](?��(?7�&?�_<�Q�?                   �       �      TREE   ����������������        X�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             HEAP    X              @�              vars           H                                                                                 ��      `       TREE    ����������������                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                        HEAP    X               �                     P                                                                       SNOD         ��             ��      ��                                                                                                                                                                                                                                                                                                    ��      ��       @         name                            	   �                           (�      H�      TREE   ����������������        ��                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             HEAP    X              h�              vars           H                                                                                 ��      `       TREE   ����������������        8�                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                             HEAP    X              (�              0       1              @                                                       SNOD         ��             ��      �                                                                                                                                                                                                                                                                                                    ��      �       @         name                               �                      (          @               @                                                    8�                      x                                                                                                                             _Ϫ>���j$?�i�I��>v�*?eB?�@y���>�|�>�-&�>��$?�4i'��T?��׫�k�>���>�%{>�t�-�n'ɋ?4��>�-�>Y�>e<�^�>�� ?�E&?���'��>_�>g{.5�?H�JT��>���>���>Dl���>�u>���h�>�*�>4Q��@9��Τ>���jwo>"�0?�</?��.K|�"�>�+?�Tf>ɽ�>���q>���>��>���0?a�_���
����£v�|��_�DD���	&_���=`1�Nz�bvㆲ_����zy.O{M1#�&�#ԯ6�/�ZW���J��ˎ���$���ˇR�̇����U6F���t�	?�	�>������?�+K>*� ?.�tV>|�>�Qd�?��
?�`������?GM�)���>��>ڦ?vJ��ۇr�e>o<�>4F�>��>�.݇�r�>���>�?x�%��>��#?e?��5�>�����'�>8!�>8?�]��>�q>��~�~n>Q�?l�?abw�X̣>:�Z�ݨ�>e�?X?�5/�5���?=�>G�>df�>�����>c��>�\�>�!�T��>$7�h��F%1�g��UQ�5<���N#ԇ�C~��I,~д�ip�*��7�.��ދ��F��l�N��~c�)���f<��-��;�C&��򆃞��2]�V�2�L�?;��'g�> ���?��>�7?��ݹ>o�d>N%�� ?L�>\'	ؕ��`L"?�)���>	�>I��>\X��`͖q��>���>U�>��?s�����?���>|��>���k�?9��@�����i��ҳ����0�`��v9��QVr2E��'��.���>��$ۆ�3"�⮍Q*�(��U�K�VD$����j���F�����jp�>�:��h���#?=.�or�>�BB���>�,�>�U�>�C�>K�>$�3;?,W�>|Ud�u�I9�>��^��?�>�?��>���@lwb`?c�?�ۗ>��d>�.��>�$?H�?����>��}>Ç��>�U#P�>�"?�F�>zY�z 
?��>R��J��>��!?�;�����?m4�\��>x8�>�P�>a�)�kQ��>��?G/�>u��>�����%?Z�>E�>����?��XA�臠���#���!��0d��������+��@��@`�{!	�l��y�������;E���1)�;�������,�R�(��	}Z߇����y�D��.�.���y&�>6B��3�>����S�?��>Ԩ?c8^?��B>f��>��?,�-�v.L>���(��}>m??uȘ>�����}�`��>�<?Y��>��?cr����>er>��>pO�	��>5<�*���H�����U��/�h1�
R;��>�>ځ���a����`���\�J���.\�-���bX�D�d?
��p��� ����Fܲ��q3��GF�=^d�̥]��������$��'��j:e���o����
9|���o8��c�b� xy[p"�chA��A@�5�H#��x/�ه����xd����7�&�?އV\Ç���1�t���X��� �b)I�>�����>��^��K>��?Z?Ϣ5?�'>�O�?�_�>h�����fA�>���,a�>+�	?}X"?��i�j���}X>�#�>��D>+��>�{�E��>w�?U� ?Pj��>|�>g60��G?(G�W��>t?��?D���Q ?U��>��և\.�>-�?9���`��7?�}���z>�ݎ>�?�P�dn��=?��>�j�>B��>� ��>B�?�N�>7� ���>��?]���,?rE{��?�	?���>kh��|�>��>��W	�>I?��4^���>�S�*��>_��>[?_�$�fڂ����>o�?�W�>��>ǟ�w+�>ɿ�>��>Ǘ���>Y�m>�h���>a����
?8
&?���>Lq��>c�Z>3h�I��>���>���o���>uP���5?���>�	?�^ŭW��E�>�2?R��>�E?AF�s��>��>J��>����C?�4?~�/���?��&1^?���>6��>w��?90�>%~��}�>a�#?o'����?��4�3)?�8$?�,?d���壇+}�>C?{(�>4�?P�����>��?� ?$���w?�o�>��⇙�?�#k	�>*$�>
�>��$�
?��>p萄�e?7�?7xH-����>�
���>1�g>='?���ꤾ���>J�?���>��>�͇y	�>CP�>I��>*z�hb?�>�>d������>����>J�?Og�>��0	 �>�̥>]0t�?��?]��P<��$�>����>]��>�m?��̩�]����>���>�Z�>e� ?����_?���>z��>?˞�=��>�o�>�p��>����P�>��1>�Xv>�M�rr?���>Q 7s��>4?d	6��A�2>����7�>m�>[=? �ˮ��R���>,0>�AE>��>D���)�>��>y�>(һk��>�gk>[��xn>_e���?>��?{q�>oWӆ*|>�NL>=lM���
?9��>ƌ5˱�r� ?KdH����>��?�h?NM /���;�>41?�˯>���>�k�켝>�c>�� ?%= 
�?�?�>���%�>�ߢ��p�> �u>�L?6�~�?�vg>\���et?�
?^#W�gć?�4��?w�?� ?,�/��3r>Z_�>Ks�>��?jٶL�G>��>��?g��5�>�=(�Ȱ06�V-��C2 Z�)<AZ��F��,�k!t9Jo!��.^wc^D���c��I��0?:L��ãb釻"&F���;φZ��h�D����P�i,�"`�������?�(�����>q��Y��>���>���>/�����>	�>��Ȅ��>��?.-����s?z��"?W �>�?7�$���W�>QU	?;�s>i'?jÔ�C�>@��>I}�>>},�&�>cb������r0	����P�1���˕Y�3�����lz��;��
���c���'7��.ڑ�*�~�@�ϴ�¡ʇ�a��Ʒ	�I�]�ч�uw�b���{軛�Ž���>���Zf�>Z_���E?���>v��>�$���>�>KH�e��>�?o��1d��:�>��%ѧ?��>f��>���������>�?
�>yE�>듒�g�?���>�d?�*0�>?A$l>������>i �P��>EJ>�.�>S��f|?���=6�K��?���>����ō�>X*!��>
�?
�>fw�.�\����>�c�> c�>�%?U9���K>$�>N��>_���"?�?íƇR� ?s����>i��>[v�>М!��>AO�>P;���>D�
?��K�?��\�{z�>��>�G"?M��������>���>��>��>#"�L�>$�?��>��.bH�>e,+�<h���@*:˱·���,+߇JK��|�,���/��U���sA���������Ňz�#+g�q�ʆ��������'� ������4.�/""����i�������]?*�#�?�)�a��>`T>�]�>^]LR�>k_�>��?�@�> �2Id���'?��w+Ȳ?5��>F��>�9�/h!�E?%��>YY>���>�� �;݃>�qn>�-�>��;�?k�̽�	����_�&�[̽�����F��l�U䪾��]��$8D
���	 ��G%�ʦ������;�tӽ\���V� �χ�j���򼽡,N����)��Vq �����ǽ�cMT�K?E���!?�Ed���>�	�>fB?���$	?3ҍ>a@�)�>�:�>��V@(;��2�>��(U�>" ?���>}�o�  �.�m>� ?J�>�Z�>����?K�>H�?��u?��>�����>8m��>�6?B7?/��g?YM;>��K���>@��>��d�5�0?�ز*^��>��>گ�>�ԯx͚�>|�>	 �>C-�>��>�����>�m?�W�>��g?���>?ݱ8>�>���?���>҈�>[��Ծ�>���>�-��a�>B��>�R��>�z�>̂H$B�?R?^��>I~����P�<�>U�?)�>��?!�����>��?	�?�p+4??�y[������%Jf$
^�`�ɏ�`
�A��Q҇���������ރ p��j���K�v�����/=U����P*���l¬���6nw�LH�����³�5��
Ƀ�g�>?\'�y�>=��o�>q��>��}>����8�>�F>\/��FE>:�?A�	��6���>Wb��R�>�6?O��>��D/bd���
?\	?��9>6$?>���ni>�ݸ>ҩ?�4�+�>Ԣ�>tkH;"?�&�?���>*��>W��S�>�zW>.6���>�W�>�WH��?�	*� ?.��>9�>8�j/�#�?�"?xZV>��>��އܲ�>�n�>��>!m �
?f!
?��߇���>zxʆ�:�>���>C?�o�3>�>�cw>����3�>u�!?�ש,q·��?䮄�^N�>te�>��><s1�]얆�z�>�?���>��?H��6?}2?��>M]x=�>n�>N�$��>x�[?x�?��l>�+�
h�>��0>���X�>H	�>����ćQ�k>�G� }>G�?%��>=ҟ�6h���?��?kN�>jC�>V~m���!?���>�Z>j:�q�>�>���h��>a��<��>a�>4��>���Ǭ>m�>�5��E?��>Cա������?w�+��4�>�X? 	?���*it'y�>���>g�>���>�-�3 ?/�?��>�]&�D?�Z?�8�j�?���:z>ܲ�>f�?ď���
n>�EF>&�"E�?nd'?
mۆZ��>\�'8�>-�?M�?�e�'�H�>#R�>��b>=��>�A���>v�>{�$?���?� �>#�Ňe
 ?*��9?wx�>* ?�d���?���>��ꇾ��>���>io4_ć?��>�4����>w��>R?h��|�w��>5�?	�?�5?i�L�y� ?ך ?^�?4���>�d�>H�/Y�x>��)6E�>#��>���>S�$���>�W;>Ir
|ő>��F>��WЇ�
?�H�'*�>�b?�
?�C;�wB��H�>�i ?ƾ�>�I?����>?�?�J�um�>�?�-��?�߆#�>�\?<w�>o̐��p>V�5>�`�>s�>>�_��q`�>V��6�>�8�>�|#?��>/�{�M��>
6|>_�>��K>5v���w"?ZcT>�i?���� ?�?b���0�?7y��>/�t>�P�>�>���>�w^>���*?x��>]ޡ��Ӈ��?�u��t�>�
�>䙥>����&�p1�>N�?���>? ?�P��/�?W�>���>B*�?z����P������)l̆X����7���?��1���4��}�߆f�C���"�ɆF��2���=+����]�������WAuu�<�>��;1�Ɏ`�Iϩ%#+o$�e؇0�_�����zmއo���
��	�0w�h=.�ėd�>��';�(4R�f#������[^�����Շ�ч0����C��G���j������$V�?!�7�xy�_��z�B�A�#�;��>�����,?������>�&�>�}�>Λ���>:7�>ZL��`�>\�!?{�p��?n�ū���>���>���>[)���hi�>��	?���>���>��ćs_�>	W?���>��̜?E�?����>�q�U�>0�?�%?(�U ?ʜ>٬
����>]�>˸����	?�4�)f��>	8�>��?=1����-�Z>��?<.�>�g�>!���q�>�>�k�>Jj��>j�>���T �>c�"��>���>k"�>�� h��>�[D>�� ?%@�>�k������>�j{��n�>A;�> �>��/+@h��>v��>���>?v!?P�?��]"?5˴>2B$?�V�b�?ht?��҇n�>���d�>_�>�N?�-�9?Kӌ>>,���>�L�>o�M�Y	�bm�>�ж�^�?�V�>3�?���*���(:�>��>���>�/?�ٞ�>?�B�>+%?D��!��>��>��:���>ӸItx�>}��>hg?�i>?d�>\D,�?��>�
�l���W�?��#��x?3�-?�K�>��-@�~%�>?/k�>�y�>UM���m?�6?5�>�?쓈>pz�>�%��`?����?�n?e�?�u??l^�>�����?3��>R.��'��Y?h���Q�>��>��?��+d0���?��>���>��>?����>L�?wM�>�$�=�>��?M���n]>C�ƅ�>J�r>f�`>BK���>���>j�x9.�>W�?�&����u%?li�)c��>�z�>^!?�`0�" f?��>6�>�[�>1�
�2=�>�U�>0��>����?{��>̽�]��>$�P?̣>]��>��>~��� ?��g>Ӡ�{�>�p�>Ɂ����pT?#�z��T�>���>���>B����t���?�Ҳ>|��>8��>&�c��>��m>�W?��	��>����J@�ܽ9�����������M\�ފ�
p��S��h�o2�����²��c�4ҽ>vE�*��+I����ݽ�H/��۫�0����`V'����D)������ f���������> �l-�>j�fa	?w�>� ]>
XS{�>��E>o�w�U?"z?���o��?sy��O�>�?�S ?khή�ǏA;�>��?���>�T
?MN���?z�s>�~�>3Q��>Λ>�H�$� ?��"e��>�/ ?jy�>|��>��>��9��?�{?C��k)�ؔ'?�B,w�}>U��>u��>(�3�YD�J�>�0�>��\>8��>"�-#�>��#?��>�/A�?ۮ�>K�}}�>���,�}>6��>eS�>��35�>��>R����>��>�}/�����	?p���8S?N?�"?7�<.B�H���>��>��>�3/?���P)
?���>��>���"?���>�����>@�`�֖�>t�?���>��Z��?�^>��,~�?̭ ?ZJ���{�q�?�闧ޖ�>c��>�1"?i=�-����8m>7�?݈�>���>�|��?���>�e�>�-"�>H	����4�Y�?6���4�������Z*w�I��$��������`,�4v�Vjه�: �M4ɇĠjL�3N����� .�Q@t��2r���/�8Ԇж	�����4K�o?5z����>��}�?�t?�>��k?l�N>�zچ��>3��>0�2���W#?��*}��>`�(?�-?��.����>�Զ>O�>uQ%?����?�,?���>�0&�>SNOD         (�                                     ��                                                                                                                                                                                                                                                                                                                                                          �      �               �                                                                                                                                             %��?���[D�?�����y�?H��?���?ז漐��?�e�?۔�%�?�p�?�"ۼ_�$��G�?���f�?���?�M�?������a�?C0�?��?��?2� 1�?}u�?al�?�@T�5��?                  8     X     TREE   ����������������        �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            HEAP    X              x             vars           H                                                                                 �     `       TREE   ����������������        �	                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            HEAP    X              8             0       1              @                                                       SNOD         �            �                                                                                                                                                                                                                                                                                                        �           @         name                               �                      (                                                                             H	     �               x                                                                                                                             գ+?���R�Y?�%��t+?�T@?��?I:5��#?R�>�s����?�)o?�1��B�)��8`?�\���/?j?-�P?۹�������?u|$?OO�>jJ??%4Q�F�o?T�b?�(?����Q�8?SNOD         8                                                                                                                                                                                                                                                                                                                                                                                                                �                                                                                                                                             c&�?                  L     l     TREE   ����������������        �                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                            HEAP    X              �             vars           H                                                                                 �     `       TREE   ����������������        d     `       �             �K     P                                                                                                                                                                                                                                                                                                                                                                                                                                                                                       HEAP    �       �       0K                                                                                             SNOD         �                 ,                                                                                                                                                                                                                                                                                                        ,      @         name                               �                                              @                    \                    �                                                                                                                                                                     |.      SNOD         L                                    �                             X       8O                             `       Hp                                                                                                                                                                                                                                                           �                    �                                                                                                                                                             o�:             (          
       �       
       �                                            �                    x                                                                                                                             u������=0Q>.m�D���{��@��>��A]�?���\"��w��n��?��?�u���>�q�?C��@��%@0���(�8�X��9��
0�Clȿ{��@fX>|�F�n��Q�@r�W����w�n�1�����£�@@x`>��v?l����rr�w,? C_����X�ٿ�F�=��@�}>r���Oܰ?H��>Ơ����z?�9��L��@vD�``��b��d��΃9�V��*�E��@O�}2�@�?�M�U!�� ~λֿ>�C��!�>�4W����� >���\@�Gh>�s�@ќ����>wN�@tp��R�ؿ�e�?w���$�AP3ŽD���`HҾ��*@�������� �H39�����@1ex��1!?�7?�"�(I�>�"��L�7?�Zy���Y��xͿ6C�@@u���ǃ�������43�6`��,�p@��u?�Ñ���ɿ��������N�ĶbA�8�@@�=b䰿��>&7c� ���^�ʾ�c>��?|")?�^#��@@�>���@�-�>�Zv���@����-?0Z? � �,z7>��5?�@虴@ er>��K>��BȒy���>���&�p �=��<����>�@��ݽ"1�����>� ?z���n��]�@��>��>."о@{�>v��>�cv=�+>���p�>���?����0��=;X?���>�i�������=�!\�^D�@@��<�?tD�� Lw>��/�(�i�8��`fJ��B0@\��?�{>@����x�>LNi� �л�N�=W>�U�=kp ?&�@���>2�;@@�H��@�>�K�@(��	^?��O���I@`�K�~)A�'!=)f�>��>i��@pn�r�9�DpR�Z��> ��ޕ�@����S�>h�?�ׯ����>�����? �-���=FN���z�@�=���,>��>�����ӷ=��ý �*@�%h?`���&پ��>?�����>Y�@��@��	>0e�_� �Y��R��𒿠g��\���5���Mq�@P_��ѿ�@��=[��5��N�[�k��>���>����Ͻ��>�@���@X�*��+�G�Z�?���P���W�����d���վ�_W�H�`���@-��Ũ��o7���n؃��ۃ"h�@�|ʾ�e޽��T�־@t�<!Q�T�@"��l�>J�v?�r.�~۾�m�>p���U���7�4|���@S� �Z@�� ��6�=�����ڥ���jf��W?�{�0�p�?Q�u?���:���B����������þ��a�`ۮ<�n�@�0��>@�+�TǠ�˗�@:��L�¾�����@O���0(A�b���+e<X�n�@��c�)�B օ�d���2Lm�xg�?�߄0���>X��X¾�3y��׽�.Z�Hr*�j���o@y�/�RS��.����G0�q��ab?th?�䅿�����+P=@ �������@H%�@��u�i��+8��m7��<2����f:�>z��?6�0?�����&@�*�=�?@��1?"9��>�Ǣ�> q_�v'�>h/[>��>�~(@-�@PK:�`f�<0�փ���`2��P�3d�H />�����͊K@����������<?���V���A�h�? r�< ��=��Ӿ�=	���L?�Ծ(���>��������[?������W?`?���>�TA����>	��E�R@�쾰�A��v����2>d�q�Hir�L4�`܀���`@���>,�n� �����<B������ ��=��D�pYl>�	���?�����\@&E� ��1�?�g>��$����v�?��߾�:�@��>��彶o���q�?�>��1��K�V+�>���=pC#?cZ����=0�p=��H�@(e=A� �>Nw������� ��?�%�=��J<P{�PO��hN��_׾�@<�.>"�������ڟ�L�R��ɾ�}�@��@�|Ҽ��!��y�=\a����>�Z��H����h���%��)^?�5����>:]��ſ;�&6P��ξ�� �� ���RE>�#�=@���j<�g�<t��&�۾������s�KWYȾ��������=�-3���~�i�'>������*�ch>)r��2u>9�%����lR�=�g�"n��|�9̓<Ãռ触<��ڼ{
�4Z�r ׾L|��f���T��=���IY�����`�=���\ ��!��!@ �}��=|�;�Y����L��ҾG���U���BA�j0��z�8޾��:�|��?�������?1T�R� ���g����$��eT ����?�,��[�о2I�������@e������/��J� � ������W"�=oǾ ���o�ʾ�I>>�w��#�s�t<����j,*�m��ɾ@W�=���x��>���=W� �;�:��'�5��C��?�������M�!��4Ѽ��쾥P��~�@�Xҿ↳�� ���6�?m�P���?+�0��}<�)�p �[�%��:��3��K�0��4��@�D?��0�GR��c�\k�dY��6�������QԨL�G��E����>L;�<���z�]��d����������?J�5��l2��Ԓ��+������/�*�	���4��uv��RD��qݾ<l��*j�����6�Y��/���x`�V�%�A:H�8`���R�F�B��)��Mm^���{�a���Bz��(mp�P.R�}0>�ˍ��ބ ����,��:�B�,�U�Q]r� ����Y�>a����}E���^>־j�����'��]�ſ)գ��p
@y�׾r�(�T�9��U4�X�n�#��m~��~��������Q�����ɉ���m�<�:��;���>��S��H���t���U��]�>�����/�m&C�n��&졿����+��`���	���h���.<c��5v��@ꤍ��wG��ԝ�����`n��}�sgx�Z���?�%l�P����@$�
�R�e@�E�z��H�ݿ����C�
׷�V����q�l��3�@��@x�S�V&���즄`�0�N��/�m��4�a����_�� c�@s���Ͽ?}w�`�?�6N���r�=�9n��?
P �0B��5V���m����?L@/�T�J�(=�sw(�� �?�D�Ė��K�@���������%�l	˾����屾ȗ��,�.�XF\���������p�i�9�q�1��WP@�e���aR����Z� ���p���1��6���t��]���}�8�$̳@��H���@��>����=�1@�C��^]��]i�j�@N�n��EA���a��,��Ϫ?�V<��=.��zD�8-�e��� �����Oc��@���J!�*$��[W����=;4�Hg3��@���׾������ z��?%���Կ�<c���@h��MB������bd�<��������d@NR�@�EJ�M�h�G���S')�������>(�^����@��?G��5�@�7?�I�?�^��#.�Z��?O��H�?�G@ �>�
x?�|+@O�3@���@�I?S;�?��\y�?�v�?���=�*��D�z?��p>�'x�hTo@���?S��>��_@ �=�j �p|���`@�%8?~�c@P;�>x:���)@���x�>(<�>'�>g�X@Q.@A �?� @hg3?�@���>��?t��>�+��P]?�$�? �;p�j>���x��> �>hC>�A��@`\y>�@#�^�g?X)?���N� @Ȩ�>�z�?0�� @HO?Dx�@5;�?�]$?u%s@�?���p�ѭ�>��E>U��@���?�w?���>c�"@И�=&l��/�>�4@4�@����S=9�L�?a�@SՖ?�H?�#�=�#@r?�?�#>6 �?r҉?�Y@?�}�>�4>3�J@P	�> @ �@`�C?0�>�?�ǁ=`哽k*<A ��@@w�=�閽�@��O> ?z:� ��<s,D@sh�?]fz��/�@
�ǿ�!�@ ᭼��,F���v@F&=v�L�������(Y.?dX�@�rI@q4� �~��O��̿s	��/���7��<ɿ��-��"�
S@�ᪿ��'�ަ@��@�H�]����4>@�޿r��?�-��2�.�?0����!�J�3�o��.<=@J��o�C�? �.��\�?ܰ��G�>M2%�ⵗ@8M�g�.'����Ƃ��C�ڌ�^���!AH]1@N�7�;��V���V�F�4L��0U�({��zn���&� F]@l_��a�@<6���ʿh@�������h�q�@o�N���(A6�o�#�PB˿���@�h�@r���Ɋ>ݙ�?tC��:.���p7��O��:n�����(�_ռ��o2��@H�$@��迴T=��� ��<
?�<����@� �̇D��qf�\�-��
��v�<��"Ah��@`� ���H��0�=h9+�h�þ�,?ֱ�>(�?���>f�,>�+@4M;>�@�@�9M?޹�4��?y6g�6A?�>$�1?��o>Z�m?D�>rX��S?�E�>"탌sm>�?�g�>�z��D�>�i�?R�?���?T�>��?w_?� :>�-�>Ir'�@��1?!�)?��?�h?�w?aZ)>���?S?��?�r�<�
�>9��=�0x?�_?p�?0�'?5q�>�.?�:����>��?8T�>�F@?6�y>^�X?X]�����>�M@��>ڠ�>�o��A�>�@���>�B�>�\��c�]?�}>�D�?/H�?K�@|�&?:1�>b�?\t�>!d�?�`���T3@?7�@k?�>@=<D?�Zk@��~>�A��c>4l�:A�=��F@Φ���B?O&?>��?Q_?\�;?i�?��P?$[F?�c�>ɯ4��>Q�O?��?|0*?bS^>�"g?Ե@x�?�e9?,�+?�2�>��f>�:.?yu@[y_?5�>642?f?�v߼�_?             (          
       �       
       �                                            �,                    x                                                                                                                             I�|B��\B��}Cn3�CZ~TB�$*D�4TBa6^D"�Bٜ�./c�BN�+ �B�tVB�EBv�A���B<}QD��D&F�Bڕ�B�:�.gJ�B"�B(�zB��t,<�LB�BLo[B�8qDי.B^��B5 BC8OB��fBW�,L�WD��rBO�cB���B�(�B�,�B��B�	rBVZ�Bf�GBB#C�G�B��BcpB�?�B�0C��pB��OBZBu�}D�@BЈBO1bBPzB���A�|�B��8BWB�p0DSȿB�[&B��-��)B�RB��B�&�B��B[��BLlvB�wdD#f�B��NClr
Bjm1B�iD�jB9y�B��#-��D㇕B��:D�"BH=Bs�FB�@FD0Be7-V/�Bʔ�BCc�B�0iD3-�-�{Bv��A��]B�nvB;��B-�xB�o;B2qBNv/By�iD_�[B��B�MB�Be+�Bأ�B��C��B�S�BJ�{B��B��B��]B��HDGSFD�`YB�(gB�GB���A�aB�APy	A3�5B	 OB�
A�]C��Ay�wC��%A��,$@Ak	-���@�2A�A61�@إ!AJ�C<�C�EA�8'A�*-f�.A��1A�6A�+-xA�":A�A� \Cӭ�@�2ANB��A��A@�	-�nC?�A��AS�XA�!:A�@TA�c�@OAJ#A� A��A7W<A@�@�AɁ?Aa| Bi�A���@�3�@s�?C���@��(A��
A˽A67�@�IA!��@��A�
�B���A��@��k,R��@
�A�M�@L�8A�W0Ag�@A��A*�?C4eA��B'�@*�@a�(C��A�h�A�q,�VC{;A�%jC:��@T��@5M�@5�HC��@W��+Y�A��A�&�A��<CI�+q��@dц@@�A�#A��4A�A��@���@�@�
zCm
A;�{A&3 A��@c�AAsr4Aj�sBE��@d! AK�A� A!I�@�jA�FAC��4C1VAwEA���@B�@�jA^�;A�!A�rBBƗXB�Ag@XC�PA�}C��BAa--ufA4ȁ*@?�@�AՙA���@[x?A�c�C���C4�kA��BA�
-p�OA��QA�j9A�J�*�2A,�ZA"A=/kC���@5�PA��B�YA��/A'f�,avCJ31AMN$A�@�AϙZA�avAF�@ݕ2AA�AA-�A�}�A�`A��@�.A��aA<B��4A2�A���@�9DCJ�A6HGA��%A��5A0l�@nA?�AC�A�J�BCڌA	�@k*�,��@A	׿@I�VA^�KAQ�`A��4A�kCC���A�UB���@�-AȔ,Cp�*Asm�A:SN*3[WCd0]A��cC1k�@r9	A�A�IC�l�@�z9*��:AQ��AX�A�zMC��+��@Y��@�s At�7A�~QA�o6A�
A���@�� A�wC�!Ab�A]"A�+�@~$eAV�SA��B
X�@�@>A�(4A_g?A���@��#A�.MC�9CuA�I*A=�A�X�@W(AE;A^�A��Ao^�A�I�@��pB��@93�B��!A���,�z>A�Z&��@�E A���@1U�@ё!A��B���B�>Av�#AD�.Ex)Apu,A\�A��^-7�@q�1A{�A�g�B���@:L4AJZ�AW��@Һ	A�b�+��B��A�rAt�SA%1Ae]FA�p�@@A��A�T�@�V�A?;Acq�@pA9A���A�dA5�@��@�@�Bf��@P�#A�E	A�A~n�@%�;A�o�@. A�ИB3�@A���@1k�-���@bE�@2�@��*A�.)A��;A�TA2f�B00_A���A'<�@}�@gcB��Al�rA6��*|W�BKz7A�'�B���@
9�@d��@h�B�߫@��%-��A��|A�UAv� C��!,���@��@N�Ad�A<)/AeA���@#��@���@�ܭB��ANrAs��@bj�@��CAf�-AR�B�;�@��A�AW�Ar��@��A��B�ӊB&� A��Ao��@q�@X�A��?b��?¿�@%�@��?0	mA���?ؤ�A\��?,�,�-�?�|1)cf?��?��?x7?���?@�A)�A��?���?�+���?N��?�:�?�T�)DZ�?V�?�e�?��A1Qn?A��?���@r��?ݛ�?3�.-���AP��?lˣ?�3�?��?�m�?=A?��?���?�&�?��b@��?� ??;K�?���?4Wk@���?���?g�\?:>�A���?(��? �?Ü�?�G@?8h�?T��?'��?��sA���?��u?%�#-Uz?~�?�)B?���?�?��?R?�?�аA�X
@�g�@l�T?t�}?��WA��?��@4�7,`5�A��?�8�A^�?�u�?���?���A��V?�S�,$��?�B@S'@�)�AQE-ַb?wq!?�R�?��?���?���?T�?<A[?D�~?=��A�u�?+@�ܖ?i9n?���?e��? ��@5�Y?q��?�ҳ?sr�?�Hg?��?�AC3�A��?�I�?��?�}#?8�?�4�@�g�@�A�s�A-_x@VB��x@��hBΞ�@UU.��@L (��2@�փ@�;f@Y�@ux�@�?Bߤ�B-��@ff�@~��+��@fU�@�\�@�,ch@qq�@��}@zM�B�D@�ʪ@��UA�Fi@��@��+&�\Bsw�@C�@���@��@�.�@�@@��@�җ@Juo@Eq*A�@�@�Ȍ@�m�@e%"A\E�@oWp@S/*@�y�B g@��@�މ@o��@��@��@d�R@#�@/E5Bm��@�GB@�] -��G@�xr@n�@�|�@��@HY�@F�@��B���@{3IAU�'@)�I@~Bz��@b��@���,~�B=j�@�GjB��D@%�]@](k@?�~BU,@� �*���@n��@�`�@��B��,h�,@f� @D�@�/�@bS�@k�@��^@�w3@�L@�K�B"b�@�:�@Ci@� ;@��@Ʃ@��A�*@_�@�@$ŕ@#�3@i�@�hVB��B�P~@|�@�``@C� @�{�@�e�Bj�kB7�)C�wCXP]Bh�D�MbB�$D"ٍB�v/=ߨB��F+�V!B�OcBR\JB "B<�B�a2D�xD�V�B(Q�B�#�,r�BŘBoچB�U,[�YB�'�B�
iB��gD�7B	��BpW�B�-hBx xB�,�WdD��{B1�oB3��B��BY�B�B�l�B �B�aB��B�,�B�B�B�t�Bzc�B5�B/,^BXcB�A/D�fOB��B� |By��B�#B���B��CB��fB6��C��jBjt2B��,�5BFcB*(BXښB)��B�a�B��B�!%D��Bް�B*B0s:B�D~�uB���B5s3,f)D� �B��DM,B�rJB��VB\x&D�BG�-�BŦ�BsT�B갅D�eF.�B>��A͡lB%*�BI�B~>�BP|IB�#B��BBRgZD�mB:�B��]B�B'Bj��Bk��B�+KC��BK��B?��B�$�Bو$B��yB�[De#DL�`BLYxB�sRB��AucrB��+B NB�BM��B��B�N�C�YB���C?W6B���,bvQB>��,|��A`�B���A���An\.B���C2D�pPB��.B�=9,�BBs�AB��(B1��+۵B��CBn�B|�&Dg��A�u=Bx�NB9��A#BC�,��)D��B�,B�qB��AB��WB�z�Aj�B8&B��B��B	WMBU,�A�!B�WNB/a/B�� B�{B;m�AM2�C��BF&5B��B�8$B���A/9RB��AFtBj��C��A���ALe�.(�A]�B,өA@B�=B\�IB�f"B9��Cw�pB�[|B}ָAVj�A��C��B��_BŶ�&N�C��@B���C�A^A�Ai	Bۘ�C�ռA��*��#B��3BmZ�A\e:D�l�-<��A���A�BK)B�w<B�m%B���ARE�A(��A��Di?B5��B,�B�An�VB� EB�b�B���A��+B�V!B�6B@��A��B�"5D�b�CɶB�\Bm�B��A�-B �BOJsB9�NC�0C;)mB��GD��oB�/yD�B�$.��B���,W�(B-�yB�\B�B}.�B`�D�rDGްB��Bw�-�ǢB��Bft�B85_+|�fB(��B��tBM��D��=B�
�B���B[�aB�7�B���*�`�D���Bl�xB:@�B�T�B���B��B�چB�_�B�jjBL�C\J�B�fB�j�B��B���B�B__B��'BC!.D�WBɘB�0B��B~�B2�B�SBykoB��	DO��Br�;Bk��-O�ABjoB;@BT�B�˟BQD�B"�BB�$D��B��Cv(B��FB5D�;�B<�B�^`, �7D@�B�3AD�1B4 QB��aB6%D��!B�@7-��B;��B���B޿Dm<�,�v+B#&�A�yB�C�B0˝B�W�B��RB��(B�~BB�xiD��sBI)�B?�^B.i3B��B�֣B(�C_�#BC�B6ΈBY�B1B��B�D�d"D�_uB�=�B9�TB��A)�zB��jA�VMA@�^B��B��KA��OC�QA�.�C��zAR�M.;�A�,@&�AːQA��;A�K�@o�A��C��WC?ƙA��{A��+HÎAO�A�TiA�5�&�;MAb�A�8TAo�C�� A;��AH(�ArEAKeA�"�,�C�*YA�KOA��A��A,ƝA�A{�mA� A�[TAL��A
��A�I�@��jA�\�A�Z�A�7bA�,BA��A�2CgD?AUŇAK]A��wA���@�ȘA6A��JA�Cj��A�?A]W�,+%A�sKAK��@	��A�V�A�4�A�$pAE4CūA
��AALj"Awx6C�cA�տA�q,-�!C�,�AN�9C`3!A�v5A(DATH+CtA�Ә,R�oA;}�AwHyA�;�C;\-|�	AX��@��PAA�lAԽ�A�iA6S:Ah!ALr(AS4CY�VA�X�A��DA,EA���AI��A)�SBhx	A�tA��jA}M|Ak)A;�VA�+zC"K)C/.PA�cA�CA�y�@��TA                       �       �                                            �A                    �                                                                                                                                             h�����&����������3(
A��f�vAXkĿ����c�|��+��&fR��|k��ٿ�u���WA8j�@��HzN��n���7�������hT�@�@-���W���;�@��m�����AR�Y3S��P��E��@Gc�Ω��@���`�����h�s����������� �/�\?P%(���)� @�<�>�����>����:��lr�@Vo��F�-�����G��k�)���*B��װ�����>�E1>��_�Q����E�Ts���h�˜2�76����v�-�?�@�^��O��@X���\�P�{��@"C������4i@�I��~��AYJ�|{�=\U��b�@8��� ��Գ�y�4��@a��[�?m1�����|F��� _��9��F�ֿ��� ̚��ٳ�`T�@�r�����Il��t��Fq�����p��?|��Ǉ��z���o`�ln�9���z�_A
մ@�t$�v����*�"�y�[;�                       �       �                                             E                    �                                                                                                                                             ���BUb�B)�C
��C�\�B�oD��BB[�D���B4  />+C�u%�"�B��B/�BG�ZBk��B�۔D�ԺDqC#�B<�"/C�UCŲ�B%^-@�B�wC�B��D���Bj�CwԏC5�B���B���,�m�D���B���B��!C�C�?C��rB���B���Bq�B��tC�`
CŦmB�"�Bx�C��qCo�Bk��B�!�B
��D��B���B`�B9�B{�dB��Ca��BQ��B�aDR8CR:�BB��.�ʛB��B�nB�Cp��B�RC���B�\�D1N&C���C��B�[�Bz�VD�~�B��/Cl�+JI�D�
CӞ|D6:�B�b�B���B	ˀD��B�C,q��Bj�1C�u+C���D�?1.mU�B�FB��B���Bt�C���B�k�B�h�B���B��D�A�B%8C���B�n�B:2CaC���C�d�BY�Bx��B��B�t�B�d�BA �D�ɀDL�B���B�i�B��JB�w�B             (          �       @       �       @                                            H      �              x                                                                                                                             �S"��e��W��e������x��Z|��*uăV	�����ݙg�鷔�ke9>����}��.���Ѿ��ž�楾��j�Ѿ�eu�G�����`���Z��þ����y<����ǻP�r(���!���9�=�i��ػ��^|=��j�p�߼2�ȾI־���5��Ot0���� ���t���&੾Ϙ�SzL��[��O���a0��/޽lyǾ�����9��cG�=:���=�)�2Y��s��	Y'���>�>���Xz������z0��W��n�_�h;��P��e��L����=�vj�_ɽ�� >�E��$ҽ�D��@��<�Fv�����A=`x:=�{�&���dr��;i$J�J��=���v5$���v=�L3�H��=���=@�_��j�='o����l|��b��Ha#>|��@t{������v����t^��x^;>�����>���;�f>P�����q�2n�=���������%�dl�=������̄�̨=B��=�i=dh��=�!v=�X�#�=�EM^�=$�r=�)�j�=�.C<6q�r�0=�V=�v�=��.=�a�;�=nՓ<��M=@��=�=�"b<�=�ׄA=��_<���=�����2=�}<��B=�/%=�`9=�C}�B�=3�)=A�H=��!=H=j2�=��=��=��=:��=�uL���S�=|�Ȼ��>'�<R7�=���<m�5=l�H=$�bq_=��<��n=�j�=��T�,�=���=��D=q2Є�s=2'�<�.�h�=� ���=�,=Lh����=�܀<�m+�d.�<��<�{�<��= ����7=�(=�w;=���=t*�=�v���G�<�0���6=อ;o�=Z����w;,�A<zy�<\7u<���<p~C�^��=��I=(�v<��>=}8=���=�F=�Ih=��:=ZW<:�rfy����=����Kq�=T�=�RL=����HD�=Z�<��4�CS!=�ȧ<���<:�<��'�R�=�&�LI��Г`����c�P}Ӓ�	ҊJ�����c�B���Wp>G�9!�Ҕ����k��n,"��G���.��Ѿ'\��-վbX���<�F�oh�ݾb� �^I��gj�(�ܾ��=�{߾>l��B���<g!��-9�xf2�]D���@��Ş�t��y_��=侺b!�gH��>�����A�^2��o���1��C%�h�%��޾�<�s���)�O���ŋ�*�r��j��~�>��`=�� �r>���=�}���=�j��@�=(p=��9���=<L$�D�[�t��=;��= ��=��=�=���=XM�=���=��~=��=�gl����=�[�>�=Q$�=� �=��у�=��9�4�=�g�=X�=C�]���=`��=�u�=���=��p=�^�==޲=�3�=�l>(W�=��8]=�=��<�� >�p�=8"�=�y�=�y=�s�=5ҺO'�=��=���=6��=X��jZ�=ԡV>�+� �G�q��[������F�e�g��o����p=�����^lN>�1Gož�>���#v�֢¾�\�ܲ��������{ݽ���,_��)P_��䨽,o�� �3��S:�\u���%l=,���$�f>�΃>#b>ެ�,�����t��.��������B��Cw��iþ Gn���m��K���P>З$�$X����;��=�Ei��b��(u.��������N�־ ��� E�<�| � U<�bJ>M�&=.�'�f>-[�=����BT> �+x��=��=o���5->�W;(~���=?m�=w�>S�=d��=m�> ��=ܿ>r�=6`>�\��>�_5Z�=gu�=<�!>=�	��)�=;��>p>#�=���>O��=\��=~�>S3�=i��=n�>�%>�>��>�k�_�38u)>�ʝ=�0>���=�:>`��<`b�=�J�=�%��">���=��>om>7b�w��=ڙ�>�%'�wR+ ��;�P���ӣ� 幼37���R��	e��Y��牽��y=<a�쯳��mO>P���O��g��8�_=�k�@E�<TO=_1&>�$'�u@��A��%>@䒽l�
>�����5�!= ש�䉳=W�
>��?��
$=�R��xٷ� (�<�����U>0�Z=pB�r1�� !�*�PO�%��>���;��@>���=q@n>�m�k���I�=�XV9�M��ǽ<��=��p�[9v�!.>&!�[c��@����'B\*ۃ�R������� �$�&ls�7.F*BU��Tr��=K��Q��E��y�lKY���=���t*����
�8,���D����^�^�
��لC�zrj]X�o�L�e�G��Z���(Bp�%����c�S8ۦ���i��3�d�8�q�K_7�%����x��ޑ���`Z�=�L������kq�`�#�9� ��޿�X'�R�P�=R]g��!.���9;����>�4��Y:���ɂ�f8��b�P>��xO�Y��ݼ����
_Q�#"��X�N�p����3���a������}�3���¹��:ab� �4��RM��2��&��=���W}D���+�@�Ǆ�ç��=�᭥�.�P��ԉ�tA3�,	&�ӻH�L�)���\��]'�ֺ��D�<���xs�<V�뽐�N�}���;���iŽ�q�^J1����T���V�jɵ�Eܻ�;OD�� ��ê.�ϓJ��ŝ�y�Մ�L�h"�B<JRӄB�V���Q���J*�M�<c�����)gY1�4Q*�"���bU�扄�< �9I�Wu�-O�Ⱥ��h�n���B*�&��u�CnC���?ڍÃ��r���������U���	�`�g�x�Ms-��J�/��@$���"�eCc��Th����Po�*ܜ���u�dsf:��d�+��i$4�?��F��vh?䪫�$�鄰�=|��=ݤq��=���XX?=�ǽ&�k�X=4qz=�r:�8�q=��>�B�;`���$�f�J�K> �5�=����8@+=p�n����=�H0���=H��z�>(s>�x�ܼ��l<��=Ҽ�>���>g�̈́�	N=@�d<�\U��[�=p�i��l >��t>�~h>�?�<��>�*5����>�RJ>�!�==�[>X�>�sF�P����Ń>�:�t>��0��ȥ>�0	>�\s�r�B>z;�=���=l����@�h�`8P���08y���k���U0{$<ɛ=�I�@� @�;R����W�z_n= p6�%ӽ�#=��Խ������k���d�1�i�8��hؘ���~=� �<A��=X�>9�>h��V�>>Y�ʽ!ƽ�=����=8Q�<�H�eҼ�½TQ}�b�b2�=S��0��
���0�O<@8+=�e	��/�,;+n.>�+��k�#d[>�2 <ņ>���|�t�P�L2׽���������D��8u��r�(��P)��S�=P^>��$��}a�-����,�E��;�ʼ� ���Zn����=�1��䖽�������P*��c	�=,3����Aq= �͜��)�X���<,���.����|�ؽO>@a�Pǽp��������<˄y36��=���L>���TtL���z�B��r?���ݻ@��g�H��<�����R�>�ȴ>�9���6���y�l܋�(B� �<�b�pm�<D����֢��*I��=2*������[>���`�Ҽ� #���S= q:�`m}<��==�V�=�o��0E�]�?���=������%>­P�d� �<�i��ھ�=aA>�����=�{м���� ��D��rXV>��=xz/�0�w=��;V�:J��}�n>�@=��><sj=H�>��佱����+>��O; �H;Z��'2>�,�����)7>J}p>��>�>H�;�L��=�j��<X�-�7�;( S�� � 2:Uq�=�,� ��:�� �?���Ľ�*>4@�=�����E>��Q=��(>9���Dμ���R/>H�3�v�&>'уF>�(+=h'>�s>�Aq>
HF_m�>H$��z��Y>�@콂��>0s�=�,�=�W��X��=�[�FM�q�=�׽S0�>���<Ά=P[����  4:H��DX�>���0w��\�>�QX��u>�c>��=}�S�^��=[��=���ֶ=3�p�aօ= �f=��9�=B�������7�=�g�=�=�l�=<��=���=kJ=��=	�9=�	�=lF�"a�=��1U4=���=�ټ==߅���=ox��	1�=�(�=�|�=%�a�{�=���=N��=�)�=��P=�T�=�;o=��=�>��=y)
�W�����=U�.=.!�=6��=���=s��<AR5=1J�=II����=Mٖ=�|�=φ�=1̤K�%=��$>�{w=����r�=I��=X;��� >��g<n�=l��=���i>���;Y�脭��=K��=8l�=ζ=f��=S	>�p=?��=m��=M��=��XL��=N42�(�==�=�+�=�f�˂>�;�O�=���=�i�=y�(�
N�=v��=��t=ix�=���=tw�=�H>��	>3�>�>�F� s��/�>�nc==>(�=^f >���=��=�1�=G^N����=��=P��=�|>�V8��=�j�N!�԰\�r!�`�t�H��=��&���x���%����0aH��E>�����P�$�t�Ծ"y�����zl��<;Ⱦ��@���ս�,��k�8۝��M�,^�L ���:��b��n���/�=��,� �::�0�=��݄vz�=�٢�������ȽT�����=P�Y�S�������r����e��� |� V,��b�235����1���h�վ�7��ૢ����(U}�(��Ӯ܃$� �P���T�����"ѽ�G�̞�\���~%+�@�x�ޜS�xI�x���?�=��G�R���꽨u�FX2����(	��j�����X����s�*$�R8�:A=	�I��i�=��Ǆ4$E����=���JG��ȃ�<�n)G>��r�R��pR��f*@�4��=�֏��B}���D�l�ҽ�x��DB�J�#[J�ڱ�=0��<v���i�T�8�!���)�`�y=7���������<38/N�=T���(���]���
�����5�d�v�)�w�����;*P�e��\1�<Ɯ��6ք���>�uަK���~.I�#�F�Ġe�L���D����M��x	:b����Ԃ1�q��_<GC�\��� Sf�#����RǄ�	�o(�u��r�f�U�oJ�b�b���kzK�����-�\0�^
���s�D���;bG�gVI�wd���Hw���,G�����=��s�40u��Ly��<
�^�ɠ�|�S��wp�>��e>O>9��닾�]���š�EU��r4����E��]����<�<E�����A5���DA�����~�u�d��=�y��^Z��ڍ=�M����� �;�_���=�뀾�2��9Ž�<~����=�T���W��oj���V�"�T)Zp���yX� ��<����덽�`ƾb ����L�Z�O;�ݶ�b��_��6R&�����R�<K�=d�½�˷����f����τ.L����!f�g�:��|Մ沺��Q�=��7���,O�6��7B��P�H�\��5�`a:��y�dJ5=��ńA��d�� �B�NG�|�l=위t=Ľ��=����gϼD�%=�h���=#0��]	� ü��=�E�>��Խ��{�Н�6��o
�|a�8[b=��.���=��v��Sr��}8�)T�0��d��������)�X�"��D��[�4�=`C�<�;q�� ��Z��8XȾI��I�־6�4���������Q�u���i>���Ϝ˾��Ͻ����̾�[龹\��z/�j∾�����W��&l!�ƾBׄ|Q��9�Z|���:�O���ʇ=�J��N�Ͻ`�*<�62 N�:2��5� �D�z������q���z��r�����ྸ��9��$�����*�+�������	оL�BID��Z�����ﾠ��,�<�����o?��Q�W�h�]tG�S�h��l+���y-���i���� >�´������e��w�>�Cv�N� ���ͨ���!���r4bk�6�݀�nɁ�z���4�I��$XL�im@�j�@��˒��C�_|*;�p����ft'\��Z�-��S^���nv��m�j���:�Oi��Gq�=�ޚ#����Qn6�6�egm�b���z2��.�vҢ�7:��d���/,��yXz�=8�&�\�F�e���7Ä�0,��<���]�
z&_�E*��T>u�s��K�r�<C����
V�@e^��{��|��"���w��X���ݓ�z�;�o����컬����׈��wτP�ʽ��<J��0��<��Z>@�8��=&>���~��FνJ	��P�i=(7���ѽL`�Zbc����RHQ�M=��A��ۼ0���p�<E���Ř�`��<�+�@a�<rg�����@/��y����*;<	�=����&ل lD�y�n����\�/���Q�䄾L������A���>U�O?\���/�����~���t�0B�ק��~��lC��pXQ�8؄0>��Xw�q��I��[��f�]�xb�R��=�T� S#:�=5�4k>�6���r�Ȱ.��XW� �=&$�ɹ<�;�?�ʘ��b�x�h|A��q�uQ�P�=5B��v<ꀃ��w���ȽDݺX�s�����Y����s�.�]��q=hσ=/���+.��#׾��羬P��D�������0���U��ܕ��>,��Le��j���u�����R]˾�U-�4��������*������|����R���	q��ɾ�.�� ����=�W�����:<=��T�-�E�����IE�$��ps����ž/O�@Xྨ��:8?�8@y `���Ҽ�:�}�����TN�0}꾣��֊���n"�vB������1_��\<�7h�����+e>8��='�~�!>u�#>Y��s�>�-�
;�=o>=�%��=�y9ڦD��">�>H>�>�g�=s�>�v@>/~>~T>`��=�;>���R�=x�r�k� >�Hq=��>����
>r08<X4�=�_ >�Y�=k��>?r>���=~s,>C��=<>)�?>h�>��S>�
>r��g�<;3>�p=\<>��=e>6�2='��=O:>}~�b>�g>�8�=~^3>�?�H>���d
��m��􋾵ס�f�\�h��.�5��&����� ���a�>b���Tǔ���z���Ӿ�
����ƾ�sd�
H��
�a�����.�M���<�y��r��9�ї�b���0�%�#��֠=���[:�p��G���֚=�^��]���ԕ��>_̾�`呾Fh��mD�؋��$g$���	���d�4"˾@^h<(�\�>97����j���.��&nj:����	ܾ-ϓ����C�+E�4<��K��|"��nA�����h^�6�����񫸾�oؾ����µ��e|>A밄�O��=W���������0�����!`پ�S����y����J ��m�z�-�d�߽����֋���$�9���?�=�ّ�ʁ���@�A�`��rf=�X��
�ھh�Խ�Ӿ��Ƽ�bj�f�~��%g� Ū�l��P?UZ�����t�Z=F������þ��۾%g��4l�;���&�Ⱦd�ھc���
\�L����J�=��ō#���y{�m�t��T��V��T����n��E���H��k�=��̃���1*��3	����ȼHw��{W�s2Ͻp�d�vH<@b�<���<���S����f�g�)n�;�9@؈��B%�<5��������u���n9��<1�����G> �:�j�4��<�j7��f����s%P�}�Y�V_I�1i����D�i=rT�C�e�+��-A��?������`�g��������B�w�*����<y.>>5=�+K�H0�����ΰ��X�����Ȅ���둽��U�f,�����=�jF���@�:�M��Uq�({�^���t��P����4�r���^����m�z������A��u��落��o<p�b��_�=粿=�����*�<���X!�0��a+���� ��<Pφ���H��㽊d�5����C=6������ܘU�tߪ=����)C�O ���~�9n�=�3C��,`�'؀=�y����-��q�;;�H����h�-��zQ������_�)�_3E��񄾾h�i�K��=y-���m�)�q��x�I��:�A��^�87��jн���o�A!�~�<O��Խ�v�Hߌ���#�8�B�=H�=�it�z�ֽ�9���F�|6�$I��\J�����a��{JԽ�t��l:�mOB�mS�.4Hb���-�OVU�<�l������޼��h����%�$�m;d����l�L�����������=n^_*m��*}�P��+"9�DwO�S�.�����%����Z�z�R�0�YR,�E�]v?�9DS�&�aL/���Z�����i/�k˄��h�'.B#)���n�?!Ʉvɠ��q]q��
��򁐄
󗄤龍���W�o�i�=(lB�e�._.: ���8�U���BQ9�=B�d��Ж�E�x�c07K64�>ށ&��O���uGL:�A`���|sl%��yX,�V>w(�=�����,>2m>`MoO+>5q����=p�=e�5���=�l���@˲>v,>c�>�-�=�~%>S�.>��=�s>��=��'>e�Є���=N���>
��=� *>"�&X->dZp;�>:D	>v�="�l 	>�I&>�X�=�>
��=#�>k=(>��>�$>l>�i)N���^:>*�y=��#>%/#>��>*��=R��=n�>����
>>w>�>ֻ>�/'�\>.:>h�"�1�Z�J��/��Ug����	�L\���@�Aő��罇i�=�)K�Zn��Y�=J����B#��q~��W=���%��8�pOF= ��=����k	�������=�]�X,s=���dH½ݒ[=�3����"=�C>�'A��� >Cn�^����AX�zw:�l]�=��Q���,�FF<�9P�J=���=(ݙ��\�=��޼@��=x�<�~�T��Rg�O֘� #�:��������P ��ڃ\�&�">�;�=��=��  ��0��� �Մh6E=&�:F�T䜽���x�/�d�=|�H�H��V=�����0���=  Q� �?�(l=��S=�%N=v�	\��ƹ��>,ʤ�>+�=��b�<�}B=x�=��[=F6z><�@�rg>���׽��=pȜ<)�> {�<�R=�l��0�A��/MI�8=\ۋ�W=>�K���u=�ǚ:�	������K ;�?>�Uؽ,>$�9>��5Y3> ��d�Q���La�m��챾�(w$U���<�[�����{�F���=�0>� \��p���\7�bľ���f�׾��K�T*��0T8�����`=� ��6'��`b!��lƽ�N�� �.�`#�p�z����=*@����RD<�Y�<>/k������J�Ƚ@r�� -Ż�4��1������鍾���uۄ�V�� ƾ�ò=ڀ����n �������b���<Č���۪�& ��~�-����P�ݽ�O�=�Y��ɋ̫���r�ف$�&j���\.B����f,�JFK�\�>�ǖ��6!����<����0���F��JG��t��<���J��ȃ=Ym����ؚ��L��P3�� �y<o��K�B�N�=¡���ǼL�	>�o�Z8>$���_�����h��#c��g:=��W��+��v��ɕ�UQ�d��@���)�B�l��=o
�x�h=e��P�����o�Yg��@�o���@�0�4�ν��บ���>�Y�;���f=`���^���x^=''��l�(��� �K=qr#�L2B���<;�����`�,���x�L=���<�U�=��>�J>v
���� =M�R���0>���;-Hy>7՝��˝���V=�˧��8��p�<���{>xg�����=�=��<�Ń>\��=��=���=Xh�<�.<��
k��=P/����>@���7`=��.�أ0��;�;�ȇ����=.����S=���=�)˄d��>�E�=���`�-�m���ʼ�x 0�����>������Btξ# T����->��g�We������Ⱦ�����b�������þ�l�6���P���L� b��ǡ� d�Z�^�ž�J��?�18�Rhy=�7�����<�2n=+Wȼ�<�ԭ�`���̽ žx���͗�Z������P���T� �. ��p�]��b��c���a�����,��vS���C;�=��!�@�̏���d+^E��=�e,���:p���v����&x�7�Y��Z����2�_��r���D>���
����N �.���=���椾��k�����ΟY���G��{ ��M� ����r·�(�����ƾ�'��R�?O�2�ʻ�=֖e�p������<Ϻ�f�=�z��쥾����SC��8.��)����T�6G��:>��tDA�3P�@�ż����5��r� �U��������n�i}�:D�۽o����������Gb��|�ӽ�l���]�d����	�7i:����������**�_A�F�>�!��|#��͟�����E
����P	���5���M&	������(�\� ��訃���Y)��CǾ�"�����:�=��ݾ��<����<��E��� ;$�*���%��[��p�<�����9������I����� ��<�v��n��ⵙ�i/�7���RD�J�;������J��>[���9�����|{� ��">澨��= R���O�����7����탧o���3�����Kþ����Ҍ�>�>6�ݝ��,'�=y�Ⱦp#��5�c�rj=�������B�RǞ�`���z38�x��ჀS��e���S����n6�T�6��͔8��/���Y>�ة>zg1�����H�˾�T��  ��u/��jfG����B�^�c���Ř��R�V\��=�����@�H����T�=74�M���C���x�� �O=`���@�C����=$�*5��`�N>�}�= X��>���=e���B>?n3ĥ>~p�=�Qi�>1�'�^�u�=�t�=��=Y>�VA=�>hߐ=)!>6�=�L�=I顄Eձ=p���;�*>�h�=��$��=�m}9oJ�=բ�=�g >�-P�=`u >�~=<Y>���=d�>n>>9:�=�#�=��>�,�>����5>	��<�Y>��=��=��<��=�Ҁ=�?�:��>Y�=��=;�+>��4h�$>`���}���G���&��C��VA�^1�ŧ��z���5��k�'�F��=/�Y�8#i���	)f���=�1s�P�ɽ�/e���ؽ�᳽0�R�pI3��C<�3��7ټW�xuw�t��=��A�U=�0��~�����<��Dz��=T����W�� �ڻ�yT��[K=H�޽6�<*�2]C�:���$���{L���}=�c����w@�_���-k��W8;���w����3�"h=@9���@��.��ϛ�hP��^^��ڄΚ���7h�J�HC���^������=%��mJ��������8�"��S��&�E�p׽\�ҽ�G�(1��$�b[#��?<!�;���<%�)������?=��@���g��Y�=i���L>qAq�������=���Գ�="1>�[��ܼ�v.G��)���f�1�$ņ�O<p����ke��p��`�x�ߋO�a�_;�5�=�圾��~��qU=|22� }G�{�Q>P�d<���QC=J@�=�+e�$|*=n��\^�=�s�;fZ�~��=�Q�<�����<TEe=��X�¨�=�!ŽvD
>��=��1>7t>�(�>�w��~��=�ܹ�$�I>(�<)�v>��ڄ ��j�L=R(�=�}|<�_�=j �a[> @�78)�<��q=å=(�>&	�=���=u�>~��=���δ�Z��=�٤�)^�>j$�=2"�=����iu<tJ*=`If�x��= �û���=lƔ=j\���>�(�>xĽ��F���� �S���؄`]����3pV5=  �&�]�0�'�� �=m������ZU>�"�qܽ�H�(��\�ǽ��r<P8�`з=H3؄�m�;�	� ��<`�Ƽ�+�=�b�l�צ�<i��,�=��f>�4����=��=��c,��b���x"� i>P'?=a;�Xƭ������.Ʉ7㊄�X>�A6>x>f(�=d;`>r�L�B4�om>��W�X�2=�!����+>����}~H�*>�؋�6K��6�.����������T���J�@;����J�>%��#
=��T��L�����ͽ����H_*�$Ͻ��������D���5�:���1��Ί�Pü�D��b���&-Լ�C��^��^C�<�򽢐���Wd���e�ᓳ<Z0�Pcٽ%��i,㽕Ly<[����Y��&�S�E������Ϸ��D��2���)k=�2Ľ���J������XG������V4�22��1ǽ�S�����>n��֡p�^�}��T{�Ӧt��XT6�E��C��Ҫ�<}׽c�=�E�$>��$��=���`q���n� �\�^������J>�$����:�r��n���kVm��Z���5�:��f=���� ��V3�=!ɴ���<��a��Wv� ���*���@-<�
9�bh�D�(��*V�$��}*� �4;ؔ�t���d���ֻ����<B���*)�$��S-���$�B�����d[���>J��=�]�;�;�
����[� �����y@�n�N�T�fG��?��?�=D���d��P܌>J&�~��`�_��JO�p�� ���p+q=��f=�h9Y�r��x��=�d�@'�=.�&�J���}=��2��ݱ=r�>�����b�=�&-��5�@W<x"��:9>pr�= ���bq�<�v<߄�TJ\�>�q�=��%>���=`��>Fe$���_�L�X>��w;��C���)���(>���J�>�H�=(᫾��#x��Xv�[U$��⑾T�j��L�#[��E��@�m>�d�辈��.��FQپr���k���Ҿ�>3P�0
��Wkt�����*ھic���W���vD�i������d	�=ȩO�`��r=�P��%�c+����b�����H��<��yN��&��8|��6�\H�#��,����
��%���m��̾�K�
�^s��,�;�o������t��Ja����;��)ϊ=�,=��.���<� �<+�
�w�=x���@=a�E=~aꃀ|�=��Q�њ��b�<���<��H<B�V=7,ڼ53	=z�=��"=��=p�<B�M|=j���<&����"�<�5��<?':��U=>T4=4�=�]�U��=���<�����=�>�U�=�8�<f��=P�i=$�<3BE��p=�\�o=2�
=��<ۼ�<R�;=Ev����<*,=��<���<\G��X�=`q`=���EQ�:�5����	|�������]� yG���#߄xH��n*>�H������B���Z���q��x���C������a�b�8��S��+B�~���Ge\Kؽ��E�@�7��K�R��>f=�< ����0Q/=���t�=�`X�د���� Ţ�@��;lD�Th���s�$�m�\��>����B�]�𓓼9n���鵈����.DK��M� ���
=���V��j����� $���4>f��My�dw��6���Rm��x�i�=�o��I�1�,+^�ҽ��U=�#Є�v�k�=��=�� ν��#����ڥ,���)�-� -�U4���d��u�*c�5��p���$�����إ �`�=<P���K�=��>>v�c ]�˝�J�"���=�	� �,���j�ڢ���ýHZ���r�PX|$=�@(�D����g��H��=�ӡ��RO� h�<��9
��=�l}����<�S�=�?�!�H���h�cn��Ͼ�	�L��	ξy�����ȾB���pxZ���<X>�;�Z���A�4����þO��~������V������{$}���6�i���M"�2���̋�8����e+�Ɇ��Ђ=|��� ��D��=�11�Ћg�&c̾M�
��Je�.�۾s�@�'޽�z�Ҿ�1Ѿ�˾�{,�Z�4��9����ľ�[�8�v�ZW�E�ž����{��vsA;�t��m�����:���?����_�>��s�!��ͺ=�7�G� m�hOi�E�5���k��fD��ս�>:R��Zn�Vb'>EA��rP1�JY����BYC�`�߼΃���ܼo߃l\Q��]/�^M<����Q�<�@�OWs�B�x=^*p�+g=O�=M�UnQ>1Ƙ� ���|J��6m��V~=����żD!�ł�5����:>� =\Q�=p�<�
>�(��\�c����:2+<��ɼ�2��xn-�^p=�Ɯ@�a=�PU=#^��:c�����ɾ+�;%����!��jں�8�����@}���iE>�ʉ��̾T�Ž<j�4ž8���u��5��6L���S���E>�:l��(پ���pG�,j��4@��}kn��]��i�r=��^�:�l��=��Ȅ(k5=��վ�㷾���Hkվ��ǽ�x��V�~������Ⱦ��Q1�TG��tg�<g�U�K��1�s径�辎;h��т�a��4;�2�>e3�ȍ܂09��@�j<�FU��(��n������M�E.��m�t�6�� �b�&� X}���1>�Ia��/D���ݾ��þ�o�����0,Ҿ$��n(����?��뎃�i��Ǿ��v8��^ž�"I��^���팾NXd=>{������t=����@Y;׍��־��c���;��սI�������p��������V�ƹ��� ���b�Ĵ�\�O�����K��f_쾺����ϻ��+�ྼ��J(�`�lZ%%����=�f�9m�踾^h���@�ߓ���,Y�%���<)�D1���a0>�eЄ2������;D%��������¾��v�:�˾Ȓ^�]�&���.���P�j����:��n��^���>�>�#���t��	=
�v��i<�_>�4��m6<\��2Q�4����k���+�d�d�������h\��j:LIƄ Aa<�d��5�� GV�@~6�QŹ��\ξ��ڽ�������{���@�\���8��pP��<�I�����m��4����}���0�v��sP�zJ�ۦ�����h�@�>���J��\bŽ>,׾�R_�� ̾�b�xo��������� ����&�"���u2������?���
��х�2�=h�m���C�<��1*�=(7��� ���І�J3�����<>��N �1O�gk��B�gx��π�o�e��k�=(wL� �ui��7"þ:�(�A�9X@�~���-3���t�u� ��;=>f�:=GP�����=��=�A�"��=����
>y�=i(o���= �a:o�e��L=x�=.{�=���=�5D=�<y=�R�=^��=l��=�\�=bg�=�F>��"�<���=��=��x�v=$�2:{ov=��=��u=0愱�>��=;�=O�=���=���=	>9=>�x=V��=�\*3�2f��=ʠF=j>~��=*�=���<.ε=��l=ĵ�����=�<8=���='@�=
�愵�=���=B̌����bj=!S�=E
�0�=�\#���=Z� =,c6��4�=h�f<�u}N��;�"z=��f=�;�=����=R�6=� �=Q\<� =�א�ƍ�=A�y��
����=��=AE}��<d�C<�CK;B�y=cY=ձm��(�=�F�=f�H=�j�=p��<��=�R�=պ�=
s=���=���Qy�7��=�؇<�@>���<�1�=�����=`�r<\�K��ן=DO��u��<D��=S���i��=��Q>��1P݄i6y�֭��^>R �Xj�����v���(��Ȩd�|8>ӐĂ��ܺ@�Pؕ�iCȾ�󂾾2A��x���G���˾yn����X
���Du/���c��w�������`��2�<�����<W�g=��݄:Ҽ�=Ǿ"�澱>��C;��X���� !���������;8���%�#76:��=�ˈ��B��2�_�x����{������+��A���z;�Z������8��<>�/j�c�W��q�)NM�����D��%�F h������@w?p� �_�
x���6w�Ä	�1����4^>P��ʄ�fq�8��<Zb��p6s��K���\�3i�j[J�,���]�����sۄo#�����)`���X]��� ���;�V̚ބ��P4�S��<��!Rt�a�G�X�������P���^�"?��w=�����a��K��`1/�: [�/� ���͢>v�4��V�̗_�8�`����x����-�*{s������~ ��#�("B>ц�0C[��>Yu��?���Ⓘ�!��M��|���I�x>Ž��<k���"�:�@�v���Z���=�o��X<���6�=D1��r>�Y�>D�B/=>�◾Ԗ��X�;�wÝ�p�=\P����T��j�T�:c���g���=����M�=�U���*>��j��ý�@����%��C�=c���x�&=��軦+��ǝ=Pg�=r.��T.�r����ݾ�1c��Y�l���ؾ9�����/���~S>�ˇ��u���4�(+�&�ʾ�[��Ò�s=��������y��D���P����� {��࿾�|^��Z�ꟽ�ޅ�=
D;���ԕ�=�D;`�U=�Aھ�2��u������V��F��3þ��о��G�&��bg�p�֚���ܽ���W�Y�_Ⱦ:g���x�6�9;p�*�}���6��pz����J� ��!�=o�/���.-���+���*O���I�pR�FT�h���⃄��Z�2�>jc3隑�P8�<��������Y�t@R�x�����u��8p����Z=q	폾�6�ӂ�H���D��u��:��ܖI=�LF��k��Q�>ݛ^�L��;><��H�9�'�ɾ�B!��'��H_b���~�Yo��%/ǚn���'=�����r�5�l�����e�����G
��QD� 1������Dɽ8(3���w�@iO�z�=��
��ud�}s�����F���|���5W�t=d������\4���1=�x�0�4��iB=~5۽8��(�׼`;�=|SؽP��=��#>l �>��� �Ƹz�Ä�B>@�?=�u`>�����$���V=L�I�&�=�U"�"y>@��� �`���^�`X@�t��=0#r=�̏=����6咽�ò����)�=�������>H 
��üR���U��:#������<�>�a �x���+3;�{Ʉ�>�'>��Խ�΄�YI����5�	�<	����u�is���`CC�42>8T��(e��l�u�0`���t������p*B��ȫ�D 彸�����S����3A�����擾2���v�e�$��Zd �2�=��2�4<���]�>��"�����(���=��M4���᏾��P���c�JO_��n��8��㴄a��5�=6����I��z��� ���釾����	��9
��hnS��"��� ����L=��r/��0Δ<�ʈ�
؄$�$�P�4��d������7��$�	w�5]HK*��	�='h�h�7�����r-�I����_��e�L�A�\3��@����<<�v�R���%�҄=�H�$Ju=U���K
��G=�`���M��KݻbD���>QH��|t�x	�GE�� >"�����2@��L�u�r�Y�0G��6x��1���2��箽��:��~�"`h���� ��<�Մ��K+�`��<NTA
9�=��>`���B��SF�����7����T��2����V���:���v�߶>m��d�����=�uþ^'|�D��$�g��H���)��g��RƖ�Lƃ2u���o�u�S��4��v*V�tg/P���_,<��V���.=��}>x�(~���S��<������[Ǿ$�T�ȯ�0�E�p�4���]�X�k��3>V$⽄�B������*��Wmt�,ա�8]����ú�B�=�Y)�`�<�P=��Y�@�\6>Z �=�'�ȗ�=���=�gl����=�1p�#	>�h�=�I���>�A�;B��D�=��=de�=�>�ɸ=0�>��=� �=P��=�K�=�����>�����=M�=�^>4q�OM�=�_�:�U>Nj >��=4�Pj�>��=V��=e�=֧=�M>:>g�>�K>�>�����D���>9�=D�>y��=Q�>ݬ�=PT�=�N�=�K]�cg�=}ڼ=���=�>œ1��=X�>ֽ$��X�H�T�@�_�T��+�!��j�ϧ�Nt��=�(�>��Ȅ7i� ���&|��e��A;�:-�"�Z�슘�������x��!�j@A�s��zڼ~T]�H$x��W���i��Z=8{���^=2 >lx2l�=����Z�{��͔<��C�x7�=h���뙽`�a���B����!��|�;�w��=k��8�2=c4����6�����x=�pR��?< ��=|%��B=��#>���=B���W�=֌=`:�7>�	��=~��=ӟ���=�#d<<��g�=��z=.8{=	[�=<�F=�G >.�=�~�=�!>��M>�d4�0B
>�Mp�>���=zv!>|��x��=
ݢ<U�=oH�=̊g=��R�O3>�z>��/=o��= �=nlY>��>z">�jz=|'�=c��#�>�>.7�=r��>)X=L>��0=��=�'�=f:n>p+�;<��=^	>�EX� ,>�»�����M��C���w߾�c͇־*�^�ز!�870���꾞�G>|CR���P�̃�B7�&Z�}�����(�!b��	��B���d~ξ�"���֦羓N��?^"�d�����?=�G���Y=dl=ɇG���@�*=(��`��·�V�^��O
��v�ž0��^���GQXτ��P�������<��8�&�;���&� �C��&��Z�X��%'�lH4��c����x��~>\!̽J���Y0��>��T0����J[��}��7��ٽ~N	>�LC������=]�����g�F�J�`����x��8v�0lm� T�!������������D�PMN� )�=4�ބ� )�o�<���Ic=�*>�X��Y�:>WB���~��ؽ��p���=�
𽬾�&h ��H��Z�Y!+���5>@��4�=��g���5=�6�5������iI��@�=]G�� ��� N��o� e�<�HF>��=׌���>Wv>�x>�/�d+�=�~�=l嘄�>��+�>��Җ>$>��>��=*s>�;#>��=��	>5��=�>�����=�P���=���=�=!>4�]�(>i �:�S+>�>?�=��>�&\�=�x�=�% >�9>6�=�U%>��=��>
�=>���=�3�U�N�:�0>�ߗ=�,>�� >m*#>��r=�6�=�1
>�����j�=��>�J:>�( >8e焧�>xq'>�g�    8ʋ������Λ��Y:�<�˽N�d��n��y�$\�=�d,.�I�4J=���I�hz��롾���vE�ءz��r��lZn=��T�J�����K$=�S�8K�<�E��їq����=rJ7� �����<�F���,�=U���/Z������ZD�-58>"�H�k���,���F��B9����Ǽ��V����=�r����g<����J�w����.�h;@��p�������}��YA�ҋ�=H*�<���i�F�Ƚ����E�o`b��rC&����@��w[H�@�D�=̢�[
��R�ս�ک�Ht���}>��g�Ccƽ	�7�\���������ýҁ�\�������½0C��S}��eA=��9�|`w���+=G$���d=��
���6�6b׽*����<�0�T$l��_Ƥ�x�'=���� �D��?a��,�ͼq|Q���^;���c&��Q<��'��'��=m۰ݽb,��}J���k�܂�l��^��M�b�ՄB2R��~��C�|Q��
���v�e����;���g���X5n���V�SJ/0��5t4	[�O�MEHo<�ߊa���h�����b��2�����Z�-�ӂ�]���b�<�}-J��*����@���t����>\e�V,<��@=����-����1�S������.�����K��<��5Z%=�?E<1-����<�:=4�6�Ӹ<C�#��W=�g:���/=�9�;���hY2;�X�(��]=M����<�ȼv��;���;S<�撄J�<|�c�~걼�&�<bv<�r��yC<��K�Ö�<9�<�s�8�����A=_-@=�t���(��*�q�[��<���2�9=A�)=n �<{���Ǟ��	=zG����z=8q<�k�<��!��Χ����<`/F���<件� �<p,�z�G񲸼�f�=����8%��2^�8�e�����L���ه���;`�g�BQ���F��|�=k!��)V�H�6�N,���tp�'���"�[ފ�GR	��Ί�c$�������b���;�X�ۼ��X� ��W��H���m=�^�bĽrw�=Hw���9 =�\�����,�˽�����"8=�H��xi�bH����P�(ob�s���˻��M��K�<*�ڽ�9��o��ح��� ���H����ʥ��\���a���;���$��>�>3$��Cq>vW'>����)P>m�b�>� >>�0Y>ꓻK�`��P>HPf>�D>�;>"^>�3d>�>>�YC>c><�P>D��pg">�D��H5>�>�WX>�����8N>�7��z[>`�<>|�>%�c��*>�b?>�&>��W>z>��Z>�R>V�[>��m>�O><���$���u>{�>�j>�D>�`>Q�>��&>�}/>a���J>j=/>�6>�o>�A4d=>������%���m�^A?���>�, �����`>�fi�����:�=:�=}�5���t�m6�����WTI��~E��g��ȅ�0�潳e���J�o��T���&�Ž\-|�\�[��?��4�j�q=�kҽRg���V�<��x�{�=��x�2����X�?�?��$}��������h(��J"�8�z��p�m2��<������0��|�`f��/�Z��j���^���G�R� $i9⿄�$����=�M�<�-ׄ������hބ��/�tW�0,a�5g4��>+���O�=/��#]G��
F��oz�j�_��43��$�@ZW�n%�B���=ԍ��C��R���p(�J��?_�}Vx��7)��ͽ�;�<Iϔ���V="�S>1L[� �<F$g��z�9=������F��Jl��r÷�`�K�����-i@�H��<�t?�p� ��K��h��<",�lc��#n�e6Q���=�jL� ��;�C2=��������w�=��<�C���n*�d')�.9H,���������G�B���#���>^���$k��*<=a�,�A�L�U�8��n7��Ÿ� ���^��n[Ȅ��3���* �~�8'�P�)=���Q	�:�:=܄�g�`6�=n�h��9�=�W�O�v��18��zx��W�=4��ܩ����t~<���X^�6�z���0��=F��qr<ڤ��t����΀ϸ@�<=�?�Ĝ�0�v���]<��=�[>�)Q=˲�:�=V%�=йS�{6�=�(����=��i=�m�_�=]���Ą�Ҹ=�S�=�a�=k�=|��=��=�d=f�=4u�=�.�=]ntE�=x�/�9�P=0=��=�a�����=P>�:��=Z%�=�7�=}�˃�B�=�=�
V=�U�=�m?=�E�=ʣ�=2��=��=���=*�����m�=�J=���=B<�=bU�=`b=��|=���=����1�=��=�­=g��=�(�Os�=8m��e�����B�ƭ�!���ھB�hR��z��ёx�_þ8�Q>3�<�ڥ��m������	�@q���9Z�~Ѿ�zξ[�ξ��Մ;��w���:���T���Oƾn�4��þ^-�=����>\�|�;��_r�/����7'���{���C����ݾE�־.�*� �DǼ�
 �����������:娾�ז��a�����Ǿ���`�ɬ
�"̡�7hq�'�,̾��4�6��N�Z�ʄܶ�HCq�l�,z>�@�<P`�/���y!=g���t�^-�ໄN�_��Uބ��K�&�+�s�|+�B���XI
�y��Pc3<�G�h���6��(�����<�R$*ۀ<_�^lI�������r�����27�%~r�Z���W��Gx���4r���Z�܍�h\��-	��� �N�X�N�z�e�_]��"o��C��L�Y�X	��z&q�����֍�Ew���Y��wĲ�^z��]��ɾ�O#�ӟ���;>��gR ��M{��Q��:&޾6�پnɔ�tM����Y�W����K7��f �K�Ѿ�P�"�d���־H�C��V�S���
P�=��`�a� �=���P��<x	�b оC`X���Ҿ�������ar�ujξ.��L�n����#�j��Δ�7Vh��/w�����eVؾ�m�)b; R��I�nh��f Z�k.q��S� r(�B�ҽ`9�D<!���_��\]��\Z��w�����ǽ\eׄ���Fڳ=�Q�_ȳ��	ҽ7�����<w�p�d�w�I�ὠW��^��=΍�=��݄P�#��g�	0=����Z�=v�τ"�罜Ɨ=��5߽����I����=P�s�-�ý�̽5ٵ���>�Լ��ȼd�˽ܼ���1O�m�����^��'>Bq��$�hM�  ���ν�j=9V1��Q0,���{��&��M�-�=Hu�<���Lk��?����6�E���S_��Rt��Nc���A�;��*=��Rgs��H��ZY��輞�M��T��x������S=!
=�tg�`=��K�}_=�����\e=�ړ�Xǋ�F��<�<��i�#���I�ź9�B��=B�����7�p]a��+C�N�A=����8�<�U��p].�	������xaX�qýW�=������۸��J�"�U�nE�:`�O���`�XCԼ��7���	�,8@=T�E>K��<��Ʉ�>^�=^�/�ڴ�=�"��^�=Hc�<�����=�k�<�
��=���=C�=��l=ܖ�=+��=DU�=��=�2~<:l�=[pV�=�'�p=ޜ�<�>0CDy>�eQ<���=ђ�=���=�5�:�#>J�`=0��=�>͘=bq�=D��=��=%>�)�=�m�l-d�@5>�����x�=�==���=⍏<w,4=�'�=����W�
>R�=�%�=K&>����%>�qZ�W���G�П�i���X�X8��2�@�.�;&0Dt<�q�`qp`u�SO�W��_��[v����a��i����!?�@ V_�o��3�V�f/��c��E�'�m=��?����f��.q��z�a�J�f$������(����zN��W�N�+���p�����9�����7��8W_�H�������SX���>���e�H�K���x;2�����>м�=N��0�;�HT.���傀�H<v΄�9˽d�\����<�!�|+>�m��ȡc��=>T�s���T�V�B�PUĽ��7�p�A� 2�:���<�\b�d�"��vM(I�=�O��m>���� v��;��<���_�>�i�>cI�'��>:́�nj�гn=a皾p�>(��=�M.�4�Q���ս[�N��"Z�Km�>h(+����=��<$�o>l=~��������=���;P�Z> ���p\#=`�=V�Y�c(>9˵>��=0�y���=�]=��#+�>.:�cBM>,D.=�ǹ�l=X�=��`]43X=��:>���=��s=Z��='�>�6> E.>\�<ӫ=�5��5>    B�>Ћ}=�u�=����w�=yg��>�s>��>RT��7N>|,4=�m�o�`>��=ٻ3>n�>�r�=W�>�w'>�\�"�AWY>�k���E/>���=�JE>6*>,�V=�V=�7;:��>L1=hz�=�	�>X�N��X> ��=�M���l�Mx��b��h{儶�~��Uľ��˾�5������`>��MЖ���o��[��MԾ����fמ�KL˾�j`��a�ĂH�]�]�����<u�^<#��x˾��)�`�J�^K��n=G�w��\#��~>�IC�
���TȾ�Z���h��'žb����������^�|�
U~�㺸��W�d�ˎ������ݽ��N�����U��DM�Ԅ;�� �bӾ(�'�F�߄����= �>����v%��LW���䓽8,�����<Ἵ"AB�W�4��>p>�,�D��!6>�:J�����/��- <2��������t��=���hV��"BL� ��=瞽�a�=���� �9����<�eټ�M�="�}> `-��j>�$��:����=�t��>���� W��Ž@�-���w\�f{#>��ԻF >��~= ��=���$x�p�<���("2=��\�.�=�s�=��9�~*A>�>�/���N9����8�/����a����Ž<����G9���j[�=�\EV�K�@��R�0����O��`7��h|��"���鑽�&�O���x$.��=܄h뼺�I��/I�8D����H߀=v�A�ޔ��[�<��Jb�=c�d�&ځ�~�Ͻ�k?��a�<�ِ�p��T����+��N��� �w7=�L��JE�=օ��;���b���c���V��`W; }�:�Z���#P�d����߄� ���K3>�wS=XW��Ѽ !�:LRy�@�K<�2��������X˼��6��z�=	8_�9���<`���F� �:����p]��AU<���=V��=��Z��$+�EJw���>p4�u�e>_�[����<��\=�Ĝ= B�<�?�=�!k0�>�$�x;���>��8<Α�>lŠ=`��= s!�`S��؛q���ׄ�^�=`��mg>+��T�=H��<����D�½v ۻ�Q�>8� �<~"P>�42��Y>�R<�����ٹ������+ƾk>���aU	�+�����Sޛ���&5>1�K�����n�	�5��?��4;ξ����J�����V�𖐾6T)���&򓴾�����O��H��QbJ�ړ'�x���EO=��� o��L~.=� �z:=�ξ��8���E۾�~i�$[�������-���א�"���`Y���Ѥ��6z�t*���e��0������2���;(t�־7_��t=���v�Nݽ��#>�ȏ�̹��ȾyǾ����Y���y��j�������7�D���h>u汄�}߾(�(=��پ"�޾���R����ھb�u��౾r���*U�b�ɾ��'��1��2���F��1��x+���= �Y�@�@=3@>�䄘�=�d����X������������b�����p�����܆���,�<<��P"뽦�!��*�;����J+�Lz˽a�2�`F�З۾��?�����[t�HI�h�'�������G��r��-�e�-þ��&�>��8#�%���B���+c>(؃SR�>J3�j��8ﾐB����*���Ͼ��޾	p������7����Y��(�!���پ]�R	���zr=3}ž��׽B�=�?�4QD�vF��q/�+����
�XJ��;Ͼ�� Ѿ���y�(_���~(��[󾝔��LKo� �Z�}�׾������%�Z�:��D���O�T����;
Z��>gĎ=�>����>3�=����=#4ƂrT=z� =�j�&1�=R�9�x @̼=⥶=�`�=F��=���=�p�=*H�=Ӓ�=d��=Y��=vz��6�t=���ⵗ=$n�=O��=�q��G�=���:+��=��=&D�=�����=7Z�=�E�={��=>!A=��=d��=S��=�Y>��=�4�R��B>�Uv=$@>�_�=@.�=�^=4�m=���=�q���{�=t�=���=�G>2�ƄNz�=��>>]�	XᘾWB�����np�/p,�p,��ڙ���:��6�ta>t4�4(F��0p<m�޾�K��{Z���'F��u��`�ҽB�߽$�ɽ�ʅq�"���P�޽]�
�);�\��|�<�C����=4>����1�=K���� ����퍾@��;��r���6>��$]�[k��х�|<���s����p�pʺ<��~�R���Z�׽�o ;�.�܋v�r�`s-�[��@SZ�(�=3��@`�9P��Gp�L�4�!L���o��6��ħ����s�l�d�&�)>�b�]����҄��v�������Tf��*G�������V"�4�����<ڢ�*���nؽwEs������n�X�i�Y�=��4����:8=d�F�=����ry��<��������s������*;��2�DÒ�7Nu��;��T��X^A��}�x�ƽ|;�|ҵ�lt��^���'��̟����ὬG��ʄ�Ɣ��=�%��ck���������^���S�A������ܾ .k�ِ����S>�[��O��;����0a���$���&ƾ��p���_�������Z�`?�
 6�Noɾ�����-�Ln]��,�=�����z�օ�=s����|<,趾|{Ͼ�彖q�����j�w��⡾j�^���ᾘg`с�h|K��bS�lض�4��@��9N~�.�ҾL�����:xPнW���r����ɽ��q�hk��O>'�a�fY��&k�������,���Bge�[�ƾ �V�a]���H>6Uu�}	���&=�{��������N��̾Z�M��6��=�z��p����������.��`��^-���FY��܁=���U��մr>A�j��*<���v}Ⱦ����Nu� }��T�r��8t�K���|(��=�6R�8V~=�@��W��� �<�̓��T¾������˺��	Ͼ�M�`3&�3>���G� 0x��*��ûF8륽D1	���������ҽ�*���Y����z �=U�����s��N�����%�n7��49��d��&��p7=Á�vb��nx(3F��Q�x�=u�/{���%�=��3o�� ��;uF >�`��}'���#���޽Dw@=p���L\��	j��vݽ�P�5xⶆ���s�Zm:=���@����b{��io��c� w�;h��<��W��7���n�z^F�h"@=��)>p!���$��P����R*���8%�:}o�p����ń"�K���!>��
�襾 �|�ʎԾ{���*���L�k�拡��(�Z[@��˽�k�8�W�|�ք�ݒ��7��^��U�����'��*E=ag.����<�L�=	���e\=2�ž!���r��Aʞ�p����H�Ի:�����%7��,b������b�<Zdd���'��3� ���`�� )ݾ��)�,�H�,臽bͣ�pu[����x�@.��8r3>��=���A��=���=d-l�<'>T&����>I��=;�$\
>.��;�n�����=��=��=Ț�=$L�=�b�=@�=^~�=��=A�>C�v����=LՕ�Q�=�M�=nx=>�O&�-U�=m�;T8�=��=Vt�=�-�=>��#>O�=��=�F�={}1>��>��,>J��=�A�=v�_�c"��d>���=W�5>���=���=�A=���=k0�=&µ�W8>���=E��=@@�=����w>��>���>c?���=��I>��2�'�>J*�R��=���=)s6���>k�~=��h]�=�>q>��ü�?�=��>j>u�>�K>d=��=�o�x�>6�O>�=��>x />:��F�R>�/�<���>{~�>�I�>I���>�s&=���=(��>7#>�OF>��>��t>�*'>�i!���a��h�	�q>�*�<vak>f��=��%>
�2>���<�ӎ������>4�<} =�Ÿ>��6�fqC>�T�������ql��|����߾&�O�ƾ_/%N�����
��M�:?�B�e>��r�ݾ��X�� �` ����:�þ����ۼ��x����C��������U|A��S� �B���,��
���]�=�;ľ�� ��ɏ������u	��w�8JC�t��2�W�����׾�����׾p���e24���曾x�uy���ҽ�~�y��M���%�H�(�Y,��?^��sb��j�T�E�􃹽H�����Y[�G+�R6L�����	��������+��=�J8�>�']��쬍��N�����ؾs��ƾ�"��z��kJ	�,䐄���w��ݒ�R���-��*��=Hؾo���}��Fy�3z��%��(�i������+Pw���۾�T����4v��$s2߫� ��+��Z��O0̾e�x�R��������T��;<ez�&����:Ó�%�[��Ak>$o�����v��B��+�+�Q5�H�f�A>�,�~����A6�0�/>d����n�>��L��r�D ��:潎����ð�~���Jo�{���|�8Y��:�5���y���7�1����x���=o����>��>��� ƹ����x���$�a�|j�Z$�4��8Ջ�3���2�2�yP�r�9->R�<��F6�Tac��(=�M��K���=�l�;�{�=bN���P����g�%w���B�܁\=P׾�P�V��RԾŐ�u����*:��6��sþp��{��*>���J���"�����Jj��[Y�w����^	f����u=�c���J���6۷~��_;8aE�I%Lg����=-$ľz�p�60۽��5��31���`��ԙ��OsӾ���&��`<d�_t��䅽�����pv��u��Za�H9?��m�X^�<s���ھqZ�8k;�.��
�꾮�3�d�����(�ܽ���=�/�I?��&,k��K��6�$x��)a��������o�o�S&>�|�����`��2v¾�p��?���=x�y]���wX���Ǿ����7���ߥ�� <������^Ֆ�Ɗ!���T���B=�-*���>6�[=]h�ԧ�:K���iľ0i��A>��ޅ��to�hMU�Y0y��v����=��;���<`��ʳz���I� AP�g����޾t��N\ѻ�?���g��@΄;p�<������+>��;ό��nk�=)��=?�����=;OCl3�<��=�`(j�=h�8���\�=��=�P�=b=���=z�>K=V=X�=�==�C�=�M��yg=#'���G=ʙ"=�O�=4aӄ�t�=�i�;_�a='ze=(Ր=)sQ���=���=jP=���=.��=|��=��z=�x�=��>+��=�}#��	�T�>�'�̦�=�[m=\�=(�mNV=�=\s^�S�=�?�=���=��>�B�e��=X�G>�#�=�d��>צ>#H*�k$>����a>�>%��[>�q�;�9��	>ru>���=G>��>f�>��=�� >_.�=4P�=��\����=�%�|D�=v��=ȧ>[�<%>J��;�@>��>�v�=�튃�>�>I%�=D��=CK�=k>��>r#>�=">��>Ytń��΋+>6� =;W>hZ�=6/>���=4e�=��>׌��a�>�7�=��=I��=E�����=�Q�<����&���D���?����8LI�������������f���@X>�VJ��� �Ի�!���[��R$d��%3���|W�l_���ؾ��X6��[L��ڳ�,�ž@����!��"��ju������<�`d>G(�˕��־��Ͼ̤@�~�Ҿ�2������m� \��>����/.�r���o��>o����3;� ��*J�����t���G; Ľ��ݾ�fU� �Q�8
�Z\�8�8�oҕ���X�վ�׾����괾�(�P��ʋ�U׳�_��z�^>��0��B�0����B�Ǿ��	�혾���P�M�����L*���4���7L��5��������B��L�=��ĵ�=�����潘#�=�!H����Ҿ��i>�TAؾv#�B���Xj��"a���\ﾂ�	�{���<��ִ�������[CL�Rs����"�}��'8	����`�!^L�Ƅ����=�qQ��[&|S߽@\����� ��h�4�Z*�">P�������ýnC�=O�!���3�pp9��W�h
�Ҙ �@@����X�I�@��;���=�g���%���,o=Pi޽h�=���@�����E=@�� ��;p�X=�h���i>�/���3�0�<z�
�V��=�����5|����������c;�v.�<yn�`��=�a�`@�԰���l��.��U�����j=���~���r�=9���>�Yu�p^s�ݟ��������@�#����_�|o���7侎駄�FҾ�25>�9���ξ��\�ﾑ����1þ$�����<gZ������`b�&�����ɾ�H��u��ۈ��}�B_)�D�a=Y8��~W���������怽V���UX�um���ž����Z��<���DO�������\��ö���Z�T���Kt$��?��¾9��'-=�Eڌ���E�ݥ�"�@�EJ>�������5>�>��{�E*q�4sM��6D��io�\4�x�	��Wu�������(��=�X~z� .Z�B2����}�k����>��B;������/�<�K�I�^6���w9<#5c����<�
�y钾��]=�Tu�#X � \���_�<RC=/z�����:�p�����I�=f��l���k$%�s�F�Ǜ9��Y �<��н�%�=�䧽p�G=�Gľb����2$�j?��H���+����� G.��?:�nQ�=             (          �       @       �       @                                             �      �              x                                                                                                                             M`p?�E?���.*�??&�A?�vQ,<�P?F5,��D?�D?l�,,/:?��>�W>,-�@?Zg?$ZF?$�M?�D�?��Q?j�c?+&?j�9??T?2��.��\?��.��B?k@?jl?��/1�@?���=�?Z?�4>?b�k?��+��?<�Z?��N?Ͱ)?�%]?�]?J�?�JQ?�?5?2Ci?�Ku-y5�*�R?�I?jn@?��C?�P?6ir?��K?�b8?�=�yU?��Y?ވC?7�^?P�-�9s?j�?��a?�0qBZ?k�a?�n -Ju?#ZX,#\?��`?��,��R?:c>Z/�,��Y?÷�?n�_?<Ie?�p�?/"p?Nk�?��=?�R?\n?k�/0�o?�j8.�^?$
_?�?[��/�>Z?��=�lw?��_?ង?��#,q�3?4�x?l�s?��F?8�}?��~?M��? �r?�JS?K�?C�'-]ֲ+ujt?�Ge?V�[?�1V?�u?	�?�yl?"R?�!=x?��x?�XZ?g�?�M�-�N�?6Q>P��=gЩ/�y�=�b�=���,FC>S��,�X�=}i�=r� ,w��=WlS<(A,���=�~>���=��=�F;>R��=7�>���=�w�=��=���.Js>~�-s�=��=��>w��.��=+˺;r��=ê�=�[>�,»�=�* >*X >D�=�>n/	>9!>�2�=�K�=_�	>���-�FH,lm>gP�=���=f��==�>>��=���=��m;��=�?>�i�=��
>Ki-�>�C>y�=?$�.�/�=�+�=���,9!�=䳔+%D�=<�=�і,p�=��@<���,���=�.�=K<�=~E�=��$>�N�=�2�=��=)��=_�=jh�.�l�=���-��=�>�=�`�=��.;��=��;Դ�=�6�=���=�L�,1��=(��=�*�=V�=�S�=���=�"
>~��=9��=�p�=k��,S��)���=TP�=5�=��=I�=�	>�.�=���=�k;�]�=���=���=E��=��h-�%�=i�?i��?.�/���?���?-�+-�ޘ?���,(	�? p�?E\H,G��?�4>d:j,ᯋ?9�?ҧ�?�M�?���?�v�?q$�?�ti?���?��?��/}��?��I.	�?i�?o�?�Em/�*�?h��=�D�?MÉ?Y<�?�v,�]?$(�?�Q�?�8p?�r�?��?ps�?2�?�?�?Td�?Kw�-�X�,��?��?�c�?��?��?6�?	�?�:�?@�J=Qx�?hϛ?%ņ?چ�?�0-}3�?�+�=<�=�//��=9��=��X,���=��+���=�|�=Up�,T��=��;e�,���=S$�=��=U��=܀>���=.J�= _�=")�={f�=B,.y��=-��-�W�=���=��=_Y�.hѷ=�J3;J\�=M5�=O��=\��+oG�=��=PZ�=Ҏ�=���=(��=%y>Y��=�^�=�e�=do,��)���='��=7��=���=-E�=���=��=�ھ=���:o��=�_�=�P�=�z�=V�-Mu�=6�?m��?R&�/B�?���?Y[-Z#�?I(,aB�?1�?�g�,5ҹ?*�>�m,���?�V�?���?���?w�@���?�Z�?�+�?lR�?���?��/<C�?��.�T�?|��?�9�?fPH/���?�R�=]P�?��?3C�?4�,�ț?�|�?S��?bK�?5�?Ϋ�?H\@���?�A�?�B�?D�.d�+�(�?�D�?�r�?���?��?���?e��?0K�?萊=�{�?=�?չ�?���?�N�-���?�}'>��>��->�>{�)�f>W��,Z>��
>Gwm,��>	P%<��>,;�
>&">,�
>�>�kT>�>�n>���=e�>�E>�F�,��>�%-
x>�1> �$>��P.X� >D6�;��>�)>�+'>k��+���=I�>�>6q�=�V>��>]�<>]3>p��=��>��+~K.)��>>g�	>��>�>)j%>Z>��>��8;R> A>k'>%�>7�,N�+>�jV?�N-?�B/��*?zJ/?oS�,7�9?Տ�,�+?��.?��D,
� ?'�=�]d+�a/?ԣQ?��0?A7?RV�??�;?�N?~�?�w$?�;?��.�QC?gқ-]�)?ߌ*?w�[?�j/�%?@j=�>?��(?�Q?cH~,�?WuD?o�=?s?FI??�I?��m?{�??S�&?��K?q"-�&u)e�=?$�2?�+?��(?pC?JX?��7?O� ?)�=��C?��B?�+?�!H?�ܠ-��S?Q@�+�ZT,�N},�p*-�O+��+s��,��p){��*��+�d1,�cn,�Y+�_o+�-1->~+S�w+���+���)��)�,5�B-�u�,��+���+�|�*W�>+�.�+ݖ,��.,
;,u_I)��W-GE,��:,��,�+�?�,s�)A�F,Rs�,�{,��*�+�+nT�,��,J9�*t�+��,�W,�޹,��*`9�)�v,�
,�߳)�L�+[�-�[:+5{***�-�6+yq<,�M?V�(?u18/vc&?�$)?���,��8?$�,�},?�6,?�,(?T�=�, +=�-?*/L?��(?[g5?�!�?�1?��H?�O?�Q#?9�<?�
�.��@?l".��-?@8-?�S?�t�.�m(?��i=gE@?,?^�N?
�,5�
?F�@?e8?FQ?[#C?xA?ǡj?c:?N�#?�XK?|p
-l�Y+�:?�=0?n�'?�'?a;?SU?uO1?X"?ڈ�<Z�B?�G<?�C*?�>?@R-d]U?AjX*���*�+�/�,���(���)���+npH)!!�*t�+��+�9�+'^�)c&�+�t�+�U�*�ϒ,�>d,���,m)�,��0)А&N�)�ߞ)g��%��(��%.*�\:,=�?+z�}*^�+�x�*���*���+�@f,���)��,<3* {(پ,�w$���+��)7�.,1+�(��(K�,�?�++�f)c�+��$~L�*&�<�*O_�'],O��+��*Q,�A�+g_+�j�*�S*�ک?�1�?�u�0���?bԎ?gFQ-���?^�-���? X�?�-;��?B~9>��K-o1�?)��?!ތ?�
�?X��?-ޘ?���?��k?D��?�?z%�/i��?�,�.m��?�ߍ?#}�?��/{��?���=��?�7�?ԫ?�E-}�o?r �?�j�?��|?�@�?��?�@�?㼚?���?�7�?.6�.�� ,�/�?̳�??�?�?|�?�m�?]�?�{�?�\=���?�g�?x�?�š?36.�b�?�6`?��7?��0Q�/?�H6?�,-��C?v��,@e0?��9?>ї,�,)?�q�=ǣN,�9?�VZ?�7?�F>?�E�?��C?�AL?@|?��-?1�G?j�L/N�P?D%.��4?i2?�,]?1�u/�,?��z=/K??��4?!Z?;�,g�?��G?pG?� ?z�O?�Q?w?�4C?�U+?o\W?u��-��])9bE?h>?0%3?) 1?�+P?Q�]?��=?�9.?�H=�K?�L?��:?�L?�� .Ŀa?w��>��>O~�/��>�%�>M�&-���>c"B,U$�>D,�>�g/,~�>�[=�2&,Vk�>��>m�>l��>�m?J��>_!�>5�>�^�>�s�>A�B/?��>�g'.c��>���>vg�>p��/�.�>���<X��>듾>h��>߆�,�>h��>Ƒ�>�Ѣ>�V�>D�>S��>7Y�>�>�q�>��-�T)�X�>w3�>鄻>�ѳ>�7�>4��>ǣ�>�`�><r<j�>�B�>4͵>`��>"w-�@�>
\?�4?ޙ�/��/?��/?�n�-~eD?��O,S�.?g1?!|,��(?���=���,221?��R?�3-?̲9?���?�p<?�fP?y�?8�,?�=<?�S/�D?�p.E�.?�o-?WRU?L*`/�#)?�{=??'�)?��N?5lQ,(v?9^F?�(<?�?L?�(H?�|q?]�@?�9)?vZN?G�{-Gpz)��=?�'2?w�2?m�'?�-??keX?��7?]�&?�<=��F?�
B?��0?GN?�V�-�<X?�E�?�&�?�N/'��?�*�?���,�]�?(�g,�ב?Nϕ?���,_=�?��@>8��+���?
]�?~��?�k�?T��?!*�?Y2�?v�|?%S�?N(�?�m�.t��?N.�Ȕ?`ޕ?�g�?�G/�?Q��=��?4M�?Ѡ�?�٭+��t?�Ԫ?%E�?e��?h�?k��?)W�?���?&�?�?�?���,���*��?���?�S�?��?-��?D�?6ќ?�A�?ڶ\=>+�?t��?ܷ�?^r�?�T�-n�?8�=G�= �.+[�=���=���+���=MC'��=��=��,�K�=1Q�;�i�*�!�=ŝ�=���=+]�=�>���=JC�=�p�=ͣ�=�ݼ=�1�+5d�=#k�,��=]��=T<�=]�N-�Ĵ=Mi&;�=�i�=���=�� ,��=�-�=��=�@�=\��=�=�=m�>���=��=r>�=��*6}+���=O��=�ٸ=�Ǻ=��=,��=ҕ�=��=���:K�=��=@��=�=Wp,�'�=6|>L��=���.O��=��=B5�,6�	>�<,K>>�9�=#��+�^�=c,6<��#+���=$�>a��=��>j{I>�(>�k>�$�=~n�=E�>K�-��>0@�-<�=D$�=x>>Sj�.F=�=���;$m>	>�d>�ڑ*
��=��	>B	>[��=�J>(W>&�)>p� >�V�=��>Zl,�g*�6	>��>���=G�>Z�
>`�>>�>��=�{B;�v>��>��=Q>�J-hf>��T?�*?�q�/�-?އ-?�Ǳ,�=?���,��1?�h/?�J�+�c'?J��=�z5+"�/?ĈO?��1?��8?��?:�@?�YF?n�?��$?�):?���.t�B?l4. n/?%0?�*S?u/,]+?�{U=��;?R�(?��L?hM',?"YB?�,7?+�?�+G?\�B?R n?C�7?2{#?EK?�~�,���)��<?G�4??�,?�,?Ce??V?23?�Z"?3��<�};?K`D?�L-?��H?P�-��P?ږ? 1n?؋/F�g?��d?,v-N �?挝+�vq?�#n?j�R,��b?��>�-(�k?���?��k?�t|?��?��{?�Ǆ?�bH?Q�a?�B�?.�x.ɏ�?K�..	et?��n?�?H�/�Zh?�ȣ=��}?h�l?th�?�,W@?��?�C|?��L?�6�?�j�?TU�?�}?_4]?y��?���,,��)y��?ˍv?�i?~�n?��?j��?�Xr?�p`?��;=�C�?�E�?��q?���?��,�>�?}5<-��+�F�,	59,/oN*�)=�E+��*G@l,��i*}�{+���+Cg,���,!b+#�F-Z�t,}�%,D{j)89>*��+kJ-2q+��+�{�,f?*psk)8�,���,���,|p�,��-(޴*Ԓ�,�
+�?�+��'6q�*�C-��+v��,�מ+�@�,��(B/,���,�,.��*�od)�r�,�Y,�,�+R��)๦,�9+�,l�I*LjI+��,�J�+y	+S)�+v�,���+b�?~g?g��/��`?�`?��X-;�u?��,NH^?-�g?2u-��[?��>�#,u�b?<��?�\c?��n?'t�?�ft?�e�?CkA?P�X?7�n?�+P/se{? �Z.h�a?�nf?늋?5˔/��[?��=TZv?�^?*S�?N��+_*8?M�}?T�t?ɐC?��}?@~?ӈ�?��u?fXU?�z�?W��-q�,DBr?�no?9�d?DZ?�q?릍?��p?�Z?��*=|?j<y?5K\?��|?T-�-��?0;?PI�> �/��>�B�>r>v,�?��-�7�>@��>�,��>��=��+���>E?�o�>� ?%�@? �?e�?8��>���>�y?��	/"�	?5�-�{�>i �>'�?F�
/́�>�=|?F��>�?v�+R��>��?�D?P�>'<?Z�	?t ,?��?�j�>�g?�@�,8�{+%a	?�?���>X�>K?��?_?-��>GJ�<�6
?�V	?�>3�?x9d-�?w�?� �?��/"��?��?\�-�
�?�c�+@B�?��?0�,9р?�93>;O�+J�?�m�?r�?��?!w�?X&�??o�?�%a?��}?V��?�[9/��?��-�0�?�݅?��?1�5/�ޅ?���=�\�?���?tc�?�',q�V?ߖ?�^�?��o?���?�!�?7�?k$�?n�}?���?ޕ�,?�,ƥ�?��??�?]ӄ?���?�7�?�#�?Ό}?$4E=g��?%Ԓ?�م?�@�?��-�0�?���+4��+0$<*w[�+�0�+K��,���,v�+���(�(�,2C,���,,��,(Yb,^nc*j�,:G+���'�U�*���+���,<�*��)���'�ޔ,�Ls+��,�ߵ,�w,8�* Ȉ+_��+I�+dV�(u�q,��,'��+��'e�X(���+>d*�k�,O�*�6h*��(yL�+��	)��*$�
)khD,�w+[W'=[�+�f�)�p�*ʺ,��+��w+�ѱ,�H�+wG�(��F*nۡ&ڲ1*�M?��,?P�/��/?�.?g��,_�:?���+�0.?.s+?ր�,4&?���=.�+�!+?��J?\f.?�8?샅?}9?�F?��?w#?��6?o��.=C?�]�-Wl+?�e2?V?
�.�%&?��^=ma9?��&?�YK?��+x�
?��<?a�=?R�?�vD?�kE?�q?g�<?M� ?�M?gF-��*EI7?��/?)?,?��;?��S?��7?CW#?*_�<0�=?��??�B'?^�B?�-��Q?�ha?,�:?�80��9?��0?$\[-^�B?��,��4?o�;?un�,y /?VJ�=���,�<8?�}`?�c1?C�B?R7�?��D?�TR?o?*�,?��??2�d/��I?P{[.��9?�D9?7�b?r%m/i�2?�o=*�A?�P<?��X?�vu,��?��H?_B?/{?�(N?i�M?�Jr?{�F?-�)?�]Z?4c�-2U+x�G?��=?��;?t85?(8C?1*g?�-A?�[0?�y=��K?ƷL?*�6?�U?s�-�t]?���?��?�l/N��?乗?��0-bp�?��6,���?�ז?EC,?-�?�II>�e�,��?ܒ�?b��?�?x��?��?^�?-}?�&�?��?o� /B�?a!�.�D�?ga�?���?e)/���? ��=�T�?LK�?^��?�-�k?���?BM�?Zׄ?��?Hm�?�D�?��?P�?�)�?�l .9��+z �?���?#�?��?$��?q:�?�J�?戴?�>`=OA�?�ԧ?��?A�?�2�->H�?��^>��.>	�.�"1>خ;>v;�,sC>�u�*��/>/V3>6��,�#>VԄ<�=�,/>*X>��,>��<>�߈>�N<>O�U>2.>�b,>q8>3�'.��E>P� --0>R�,>�kW>q��."�(>E)�;�?G>��3>�V>8wV,��>��G>'&H>]>�H>x?M>lZt>YJ7>�� >n�S>3�+6��*��D>�@>�k1>�/>o�H>�$[>8�C>�*2>�\�;�=>�9I>�'5>D}T>��`,��N>��?��O?���/�W?TT?�-�qi?:c�+�S?� S?(,�E?.7>��H,+kV?��}?ʋR?v_?�Т?�b?�t?`�3?G-H?�f?ـ/(�f?:[b.;aU?&�P?�ф?�[/��K?]��=��b?�!P?j�?�`�+��,?��r?��d?�;?�^p?u?N�?D�g?��F?��y?_�-N>�+�|g?�Z?DnN?3)Q?�l?f
�?�|[?}+K?�&=v?h?=Go?�X?�m?�:o-��?��j?��@?�w�/2;?@�;?�AW-�H?b�,�oB?�8?*/�,��2?<��=R�,1�=?� h?�?=?��F?6s�?�G?��W?��?[C7?e1N?��*/�T?�	D.#U;?"�>?��l?0�/��>?f=�CN?p�<?S�Z?M�+�?�%O?l�H?�'?�9T?��U?�p�?�qG?��.?[4c?��-݀�*��Q?�B?{	;?��??p O?[�m?T�D?J;?��=/�T?F+M?�M@?��Y?�C�-U�l?2�=��=��5/���=5��=t�,~5�=�Ĥ,.��=�,�=B++I�=�o<M��,&�=���=9|�=�&�=e@!>��=��= �=���=��=��.��=P�->�=��=���=�.�q�==�;Vh�=�@�=��=M,�=���=�
�=43�=7��="u�='>���=/�=�D�=se�,�)o"�=?��=5��=(�=·�=�>���=���=�̍;Ҷ�=��=B��=AR�= -ԭ >�E�>�'�>�h�/l��>/�>�*v,A��>��L+c�>qp�>�th+�Y�>v�=�]o+��>���>�5�>;��>h?u=�>ɺ�>��>���>O�>�̸.���>:�-���>���>t��>6Q�.�-�>���<nm�>�f�>JT�>��,�K�>6��>+#�>�l�>1�>(�>�	?�{�>�V�>1��>�m-h�,���>�V�>b��>ʁ�>0�>���>:Y�>���>D�<E�>���>���>�I�>Q��-��>��?3L�>>ۼ/��>�g�>S��,XD�>uN�,��>�.�>H4,��>-l�=:Y+�o�>�	?��>_9�>�7?���>*?�V�>��>8��>兡.�n?>�.g�>rk�>O�?\2%/w�>�.=��>G��>�?���,qJ�>�t?�.�>���>��?K�?ez?�D�>�/�>��?�Z�,3Q�+u��>!%�>#Y�>�v�>	��>��?m0�>">�>��<��?��> ��>�?u�p-��?���+O��,7+�+B̆)\ �(1?+Hl�(���+cw�*�{
)o�,�g(��,�&*��+�cf)��F,B�,7�0'`��,�Ф+��,��:,� ,�&*G%,�}�)���*i�P,u�*�<�)ў�)&ũ*���)Ұ�*�z0,t�*��(f8�*Z�,�n�,�=@+�K)��,E
A+�e�,b�3,��+ ~�*)�+
&�*ё,&P+c��+�vw,��5+��,b-�,F�('P+�%k,8DC,{�,��J++8>e��=F�.�L�=0�=���+�C>��*7s�=m��=��:+8��=�!<�ǎ+���=G�>�N�=7|�=�=>��>Ώ>��=z��=��>8�.%*
>?�P-��=;�=l~>J�.B�=~z�;ʜ>5<�=c.>��,���=t>��>��=��>)�>�D+>�v>��=�f>̉+��*F�>�>t@�=X�=-�>��>��>0��=��C;��>א>���=pi>Z��,%�>`4�?��M?��/:tL?E�Q?z�,z)c?�L�+��O?;�O?k)�,i�G?3�>���+M?lqz?�P?��[? c�?!�c?��u?� 0?HG?̴^?��&/�if?��.R�L?xP?wm}?i3/R#J?e��=��_?�XN?�?y?��J,�(?��i?6�]?y�8?��h?0k?��?[�c?G?�u?�{-췛*��b?�iV?��N?wlI?��`?-B�?KsX?��B?��=�c?�$d?��O?��o?��-n�y?�_?�78?M�/p 5?��;?(�=-&�H?I9�,v5?�7?hl ,�-?���=�+�B6?\�[?�[9?�@?�R�?�GD?v�S?��?�1?�ID?X6�.*�P?X�$.=?�/7?�dd?,�2/v4?I v=�@K?W@8?�6`?�ڸ+�%?�J?��G?W�#?�fO?�tP?�z?��E?��0?JY?
I-~�=+�J?A?�t9?�@<?M�O?��^?٬>? �0?-�=��J?�O?��<?ӁR?P\-r�b?`��?�)k?(�g/��c?��k?S�_-��?�,M	i?#o?�I-�[\?`F>���+u�j?���?]
l?b�{?]P�?��z?�'�?%H?�b?~?�5/?��D.Bs?�l?���?��Y/8�g?뗛=T�?�Ll?���?��!-�@?���?+2}?�_P?X��?�.�?���?�|?��]?�.�?v7.�,,�Ȅ?u,r?�Hj?�l?� �?�0�?�Rm?�}a?��.=���?/Z�?(np?O'�?p�-��?�ؑ? o?D�0�?k?[�n?K��,�R�?��,��p?��r?��,�xh?>7̌+�ns?��?Fh?��|?���?�t?�S�?u\L??�d?�z?�:/x��?V�.Xj?X�r?��?��B/�j?f+�=`C�?��l?㨐?�Kq,�C?n��?�Q~?��R?kA�?/�?��?x�?�p^?���?��F-O�,�l�?�z?/r?Ym?U\�?9Z�?��u?��h?R+0=���?*؃?�n?\�?���-�ݍ?�/\?;'4?�ޯ/��5?Q.?�N*-�<A?C�-�4?��1?~G+� +?�6�= ��+p),?C[V?�/?<D??^��?�F=?.L?x9?�5,?��<?b�.#DF?4�Q.t3?�7?��\?�fj/�e3?p�a=��A?m68?3�X?1}�+��?^�F?�>?��?YG?(RL?�<s?�bB?��#?�R?}m�-~6�*�!A?`:;?8�5?A\1?�1B?��`?�N6?	<+?<<�<rD?M�H?�g1?7�U?���-�`V?���?�qT?�Qy/�R?Y?x�-��i?'2�,cY?�R?��l,��D?+></�,Y?��z?V�^?dpb?��?��g?�dr?c�3?BpL? Mh?;��.��t?4р.�1\?�AZ? ��?�ԅ/�gN?�Z�=$�g?.#K?�%w?�=�,�I-?.Ak?��i?��=?V�z?�aw?M�?�d?"�H?D��?�GX-@Ϯ+�Ul?�W?�U?1�V?�n?���?f?5�K?r�=��i?Mn?E�Q?b�o?S��-�	�?t|?�4Q?-$�/8pN?��N?L�,ge?��-��K?uP?kx,�'D?(>OP�,�qP?ex?\�O?��[?Sס?k9]?*{m?\2?H/G?3�`?��.�	i?��.[�S?�'U?�}?bW/6�E?�0�=�X]?�GN?8Rw?��,��#?ߎg? �b?9@:?�l?��g?�ŏ?�s`?�
H?��n?e�-���)��c?oAU?\O?j3L?Eg?VRy?��U?�7D?rd=`�a?#Gj?�/N?��g?��-��z?K2�?���?2��/�+�?���?Y�-Р?{�,ŕ?
k�?���,���?\^J>&�@-�ߑ?Њ�?g��?+��?I��?Ӳ�?>��?�w?�t�?��?��%/.x�?k�o.�?���?Hy�?��$/p��?�=���?7��?�d�?��+��g? +�?���?F~?V�?O��?�d�?�q�?D��?Z$�?G��-m�q(o�?�ט?���?\�? �?���?�(�?@��?w�^=�D�?���?��?T��?��-ݲ?@}�?�0�?��/�8�?��?��,ݜ?�Ѐ,y=�?X��?�T�,��?/;H> � ,L
�?�l�?B{�?Ɉ�?� �?�B�?�ѣ?;�o?�P�?�g�?��/�Ԣ?/;.(�?97�?A��?��M/�S�?c��=�Ԟ?KĈ?��?��+��h?���?g��?rɀ?h��?b��?HK�?_��?�Ɗ?[ͩ?P� -l�)-Ι?E�?-\�?�+�?�͟?#N�?"��?�|�?;�b=r��?J�?{��?^�?޿^-a�?Ao�>~Y�>�:>/?�>�O�>�,o��> �u,���>��>�/,�ā>g+=3e�+��>)@�>�H�>���>�,�>J��>!�>+�n>�L�>~ �>�>�.Ś>
�.�3�>�Ԉ>�\�>��3/?�>?k�<��>i��>�1�>;E4,)�j>���>�Д>oHp>�Н>Ó�>ü>��>歂>�G�>�ud,! �(�U�>���>ӂ�>��>��>�?�>Nb�>\�> �J<ib�>�&�>�W�>�i�>'�-7K�>�pp?GZC?���/,�A?�F?ާ�,J�U?oI+O�A?�QF?�T�+%�:?�[>�?>,3F?$pe?,�D?�>L?
a�?�CW?��b?B�%?ړ>?��R?���.	�Z?k��-� C?�KC?�w?qC/�e;?�׈=v�R?ۈC?8�k?ʊ+T#?�D_?�V?;�.?�b?��d?�b�?�V?��:?1l?��},ǳb++�V?�N?�??��@?�\?k�u?�O?Q�>?�� =^�]?�	V?��B?��\?�Ū-٢r?��h?�o5? 0_2?�t9?ή0-�EH?��+�8?��6?�d�,b�0?� >Y�B-H�7?��^?�k;?dA?�h�?��D?��R?DR?��6?$dM?oiK/C�Q?֑,.P<8?57?��b?��2/U�6?}��=�zI?��2?�a?h�$,��?��J?�G?�B$?[�Q?ZT?��t?�6H?Ja/?%c_?��-�y�,�EO?8�??5;?�B4?�LK?�E`?z�@?u>4?��
=�J?��M?>?�WW?��-��f?���?ɺl?."/�i?��n?��-VR�?῝+��f?��s?yVz,;�`?�>��`+�o?S��?	Tk?@�s?t��?�c?�ʈ?��J?�b?;��?�/���?�
.�Fj?D�l?��?<�/z�d?L��=0"�?Hk?J�?k�,�A?�h�?=��?��Z?��?�?YT�?-_�?��e?�Í?@gZ, �p,�?�Uy?�Gk?һj?ă�?�?a w?�]?O�?=���?�m�??�n?*�?��Q-%��?�Ú?U��?%">/J"x?;z?75"-�.�?��=,��{?n?"�+|�s?8V,>!�,�{?`��?�|s?�E�?��?"̇?���?� X?�Sv?�x�?�U/��?4�-s��?���?���?g�/��}?��=�|�?�b�?�G�?`��,0�O??�?W-�?9�d?A�?� �?�	�?'�?zVn?��?���,��	*l��?��?�Mz?zwy??��?Ġ?���?��p?`n?=�Ռ?u�?�?���?,L!-4Κ?R� >h>�/��>�� >���,�>�J�+1a>(��=��Y,N�=L(�<'��+>q >�">�a >a>�cN>�>��>��=���=��
>$�P/vb>��.
>��>�d%>d/J�>��<,>�	>�j>�"�+D��=��>:d>.��=U>��>�=1>�E
>���=��>��,��*,c#>Г>ǫ>u�>B�>��+>¿>7�> ߙ;�>�o>-�=�!>/�-AN >��:?�&?#$	/�w?�?��9-��#?�i�,�Y?�H?)Q�,>�?�u�=��+m?�:?Rr?'�"?�`l?�.#?��/?ng�>��?�#?a�x.�*?{ֶ-�M?d}?�g;?�t�.��?4�@=J�#?c?Z5?��+-5�>��*?��"?�e?��/?�j)?~M?�z'? �?�5?��e,��(>1$?� ?JE??v�&?H<?T�?B�?�5�<�!%?F�,?�?��.?8��-4�;?Z|�?%�?��/O�? ��?l�--|�?p�,��?���?z�,��?v�y>Ϻ-?�?f�?��?/��?��@�P�?�B�?;Ж?�6�?�"�?X /���?ݱ.��?$ڲ?���?���/r
�?�r>m%�?r��?p��?tަ,4ϓ?�T�?��?â?f�?���?���?6��?Q{�?ۣ�?L��-Հ,Kq�?]��?�z�?I2�?99�?
�?tz�?�C�?kp�=~��?�8�?�o�?��?�]�-6��?���?ߥ�?��l0�6�?���?�e?--��?vr�-*�?p�?$W-J��?O�_>�V@-�y�?��?%��?ά?2	�?��?_8�?���?�>�? ү?ɟ�/$��?�&�.PU�?�У?A��?I'�/��?ߡ�=�I�?g�?�{�?�Ce,!Ѓ?Z��?��?}��?���?�ӽ?��?6�?ك�?\��?ׯ�.�|�+���?�?SW�?�?�?�j�?��?xg�?�j�?%�s=���?N�?��?T?�?��.���?y"�=(r�=�Y�/dC�=�	�=6d�,��=׍D,�=n6�=�:,�:�=v<��+ �=7��=���=	��=��>���=% �=Xϗ=o2�= >�=�\ /)��=��!.p�=���=uQ�=��.Z-�=��;f��=�=�1�=���,7�=�b�=� �= �=
V�=���=�r�=/
�=_��=ג�=+��,
Y�*g^�=y��=��=}��=� �=���=���=i�=�1;딿=K9�=:�=q��=�n8-Fa�=��d?t8?�!�/UQ6?��9?��9-
iE?d�,,��5?<=?� -��/?+��=QH,n�:?��X?�8>?�D?(~�?�G?�V?+^?c�-?�OJ?��I/��O?��.�,<?�9?.ze?v1/'�4?�w=��G?�99?��V?S��+��?�<T?g�H?�$?ǮU?ǇU?n�}?��H?CE.?W^?R/-@�_,�9G?$<?׏7?� :?{�F?Za?��C?�t/?2�=I P?�tK?9	;?P�R?��-gFd?�7?��?��/	G?��?��7-�!?]x:,��?��?�~],{�	?�|�=ً,�?z�.?0d?�n ?@jl?|�?��,?2��>(�?�5"?gq/z�'?N	4.�P?o1?ߵ6?��/SI?P%E=}�!?:�? 80?ޜ,H�>��"?�J?c?��#?7.?�1N?��?�n?35?w�,p),_!?�!?uC?�?�T%?ڃ7?�?�?=��<,%?�8&?E1?l*?�	4- :?[�?/t?@�/�m?0�t?5��,oH�?	E�+տs?o�z?���,�d?�">E5�+p?�k�?�v?��?�½?8<�?}��?b7M? �h?�]�?y�C/��?�a.�	u?3fx?Ǖ?�H5/~|j?�@�=���?�j?1�?�B#,��F?�w�?�b�?�T?�?�w�?Vk�?�j�?Eb?:��?�?-��,A2�?��?[�s?7ho?�B�?�_�?��?��k?�[:=���?�Ո?�$}?Kh�?�"-*3�?�X�?�<t?S��/'�i?b�o?R��,3)�?_�,�o?�q?��F,k;h?�$>bp,	�q?�o�?�;q?\�}?�ĸ?x$�?��?��K?�md?u�?���.GD�?���-��p?��s?��?�%S/�$j?�,�=�?��l?_*�?���,I�D?h�?��?.U?�g�?q��?&�?�u�?u�a?�p�?���,0l+��?7�r?:m?w�r?q��?ko�?Ew{?Dbb?��/=��?��?ar?�W�?�Lz-��?2ʠ?�ށ?)/֩~?&��?�~-�t�?3�d,X.�?|��?�N,G�v?��'>��+{}�?+j�?ۣ�?�v�?�q�?hR�?ȯ�?�f[?b�s?��?��\/<�?�eS.��?��?� �?�{/~?�=��?q8�?�?7f%-�V?蚑?��?�(g?��?\��?���?���?�/r?M��?6.v��,���?���?:Á?@��?_��?=�?T��?H�v?��@=�͐?�?o��?f�?��H-?�y}?`iS?T��.��H?�K?�K�,��a?+2�,��O?��P?�@�+�"E?� 	>��8,n�M?6�s?� R?{\?I)�?c�Z?~Kl?9/?PC?3�_?��.�f?�h�-�]P?[�J?8��?���.�tI?v�=��\?��N?	�t?�,#$?Kg?-�_?.�2?��k?g?<T�?td?�hC?&t?d�,��{)��`?ptR?�nJ??N?yQ_?�C~?��X?�@?��=\�f?�se?��K?5l?�Xv-�Yw?U��?��?�MH0�J�?EA�?A��,DƠ?R�-��?�K�?�W�,i��?4�E>�/d-��?�?1�?�p�?�u�?0�?>�?�}|?jύ?�ס?E��/���?]�.� �?�>�?;��?��/1��?�T�=�*�?�Ŕ?�j�?$�-��p?�L�?��?4g�?�h�?<e�?U�?H_�?r�?���?�TB.��\+���?�Y�?t�?%ޔ?���?7ϼ?���? ��?��b=�Ŧ?��?�ʕ?=�?�.y�?61�?6Z?!/J�[?�
^?�-��o?vJ�,�?^?��[?��.,jLM?��>�{�+.�W?�܁?�P_?�'m? M�?8<o?T�?�9?R�T?�3r?��F/j�v?c�a.�V?jGX?-�?�I/�HW?t�=j�l?�nW?�2�?aL�+�:1?�Oq?��c?�F?��t?�x?Y�?`j?�SL?j��?i�.�,�cq?��f?�r`?7L\?��o?tr�?�c?�R?ϐ'=�Ww?8Yv?G�Z?�?J6-:��?�E>)T�=͐�.6'�=���=($�,ĝ�=��Z,��=S��=^��+���=&$H<��,�}�=��>M��=���=�*>l
�=�h�=�6�=	��=���=�.n9�=!�A.E�=L�=��>�F�.� �=�E�;��=���=?e>gz�+v�=�k�=��=S�=���=�P >>���=���=+��=ъr,;+@)���=^5�=B�=���=��=�a
>o[�=ވ�=��\;M��=���=�=�V�=g�n-��>�F�>�k>~�
0�k>��d>��'-7�y>KKD,b�g>�Ig>�,W>��=���,��`>�U�>mh_>Q�n>��>�Sv>�m�> E>�]>��o>8�/*x>9O�.�[g>��f>�@�>Wi�/_�[>)��<t�w>k�s>���>I:$,��?>`<w>h�w>�F>��>^+�>I(�>t�s>^�P>�؄>\k-C%,MM|>1�y>�h>��_>8�u>�S�>i�q>�!g>vY<��y>��{>�V>���>F�-Z��>�μ?�S�?+�/��?9͖?�n-C˥?Wr�,���?|+�?6��-*�?��R>Uؘ-�W�?�^�?D�?���?p��?�g�?�>�?���?i�?��?��/DK�?M05.��?o�?;>�?3ݗ/=v�?��=;�?�#�?	��?ڌ,O�z?��?�^�?V/�?� �?��?T��?�]�?d̎?�_�?���.��,�?��?��?^��?=.�?rپ?���?�Г?��v=�(�?
��?'g�?���?X�-���?kx�*�C,��)��,jK�,�6($�l,,,�e0,��!*��c,]��,�ָ+�Ȯ)�B�+]�-�̌,�Xo,�8'��)�?*�*a]J*�5*�o�+�8m,OwM+U�-*��F+�C,�%���*�Z�+l&#+p+�`P)|�.*���)h~K*	{�,�,+�� *Z�*;�+hx�*N��+���,,�d%(rV,3��+���*~)�)K��,p�+^e�,�.�+`�`,�8�,���+	�,��`+�=+;�,�F�?0��?zT20%��?P7�?�M�-�D�?9^,��?��?�,~��?��M>�*q,/�?�ڷ?x��?Ik�?�7�?���?���?�΃?���?�b�?���.Ю�?hHf.똙?'m�?��?�S/��?K��=��?V�?���?�-�,Nz?�,�?�.�?h��?�Q�?W}�?ڪ�?0[�?���?�?�h�-�yb,O6�?��?ߖ?�Ǘ?}�?衾?��?jH�?&�f=��?��?��?�ۮ?�-_v�?���?r��?�-04�?4?��}-Cݎ?	��,q�?��?�(�,c�{?5�)>P��,]��?�m�?�L?#��?I,�?���?
|�?�Z?˝w?�0�?�z�.�?�C�.�~?Z��?`�?ٽ�/1�~?�=M�?o�?	�?��g,�iT?�'�?V��?��b?���?;��?U��?FY�?�t?V3�?��.�r+\5�?D�?�W�?%b�??�*�?O��?cx?�n8=��?�?�~?h�?���- -�?c?��5?h�W/0�0?7?Ԇ+-�G?1�,�9?c�6?��Q,j.?<�=�>�,0=8?�eW?�	<?��B?}�?/�>?��R?��?
�-?�9F?�=�.b
L?6 .�29?�%;?g�d?$e0/ 3?l�y=i]B?��2?��]? �e,s?��O?P�J?�[#?O�S?9IO?��y?�2F?��.?�Y?��-� ,e�H?�C9?��9?�5?FK?��a?�B?��-?>=;�H?��K?[�8?THQ?NX�,'hb?���?{�L?���/CK?�iI?�e5-fg?��/,ۗP?�eO?n�2-��F?c�>�"�+�3M?R}?k:L?DV`?�?m�Y?��m?�0?�+G?��Z?#/	�j?3�Q.ɭQ?/�L?�
}?�y�/:�H?��=�c?}Q?�&u?zG�,ah)?f�f?˨Z?N%5?�uh?q�k?�?�a? �@?i�w?`-�Iv,��c?�{W?=cN?�GM?�e?�R�?�Y?sA?Ni=��d?_�e?6L?�l?*(�-r6~?>ބ?�W\?�M�.��^?��[?lsp,�j?�3-�EV?�b?l�,A�S?#�
>��,��]?vM�?�K[? �j?J��?%;m?x�?�N7?�T?�j?!3+/@p?�d�-�_?� Y?�?H7/xW?���=�9j?�$b?�z?��,��5?�s?�j?zB?��y?���?֜�?h<p?(;M?w�?׌N-<G�*��x?��g?��^?(RT?�r?�?�h?Q
T?b=�r?��u?�'\?�I{?B�V-�^�?\�`?3;2?B�K/Nz.?�22?Vύ,9F?[t�+g�0?�w0?x~+��&?�A�=��,��1?�Y?vY,?�i:?���?94??}J?��?9I(?)Q@?��.֖D?@G�- �2?�,4?�3a?�;/��.?d=�d??�93?*yR?��?,�	?�{F?�<?��?<�J?CN?�2r?'7@?�('?�T?�Y�,��E)�*A?�9?�I3?g�0?�B?�	^?-:?�&?���<6�A?x�D?�65?4�K?V�s-TV?�ޕ?(w?M%R/X�q?��t?a�,���?I�X,��r?��q?JoY+�h?CS'>s��+Qt?&\�?�x?�s�?�*�?�6�?�Y�?z�L?�Qr?F��?���.���?4�-kw?�w?��?l{�.��v?���=K�?�n?�8�?�`�+DH?iI�?Ą?�$V?�<�?S��?q��?ۘ�?��j?�ݓ?C��,ùQ)���?S�|?G"r?U�q?�Ň?Ӽ�?F��?�Ye?4�B=���?���?��y?zz�?mq�,�E�?M�>���=2�-��=���=d�+E�=lS:,F2�=m��=���*'�=i�<�+�x�=I��=�G�=l�=�>">��=�o�=�{�=���=�O�=�7-��=�I-�l�=2~�=���=�#.%��=�7z;�'�=���=qb�=��+a��=�s�=���=	�=���=J�=��>L2�=�h�=r��=D��+eN�,��=��=Ku�=���=�$�=a��=��=1�=��3;�S�=x�="��=�m�=1�6,���=6�?a�Y?j�/3�T?$�W?  �,an?�5�+�W?��\?�M,�O?��>��,��U?'�?�AT?1>d?��?�?h?��z?��6?��K?��l?L|//&p?��-%Z?/�Z?�څ?�N /IS?Yɓ=�f?��W?:|?�l{+�+?i]q?��i??r>?�cx?��v?�?W�k?6fO?C/�?��,
��(>�m?X,Z?�PW?)�P?�o?]��?��a?��P?��%=rm?{�t?�bW?us?�"$-��?S�2>.>�`�/�3>�>�,�,��>�?�+�/>g>�s,�4>���<��u,O�>l�(>!�>��>#�`>�>-#>T��=��	>k>�7/��>X�.�
>��	>M�+>�`/��>T�<�)>�`>�Y#>�:,`��=a�>�>��=7~>#J>Ŀ9>��>w�>k�&>wg�,�A,�[>�Y>��>p>��>v$2>��>Fk>���;:�>->�>�T%>��-+Y(>���?��?4�/|�?f��?�WX-C�?�3�,�M�?�8�?�״,[��?�]\>�[<-Zȡ?>h�?=�?rh�?��?2�?��?]��?�'�?�
�?M�</06�?�s�.��?0̟?���?ⓑ/�
�?�<�=d�?y1�?��?\j,g(�?!�?T��?l�?b��?��?F��?��?�^�?�7�?�.�{�,߬?2�?Ko�?'_�?�?<��?�?w��?�um=���?Ɇ�?:�?�<�?�-J�?eΘ?Dx?�D�/�5z?�@}?C�,��?��8,�|?+1}?�ǽ+�p?�%%>�|�+	�x?�S�?��{?�j�?3�?�؅?�Ύ?o�U?I�r?fm�?��/���?-� .�~w?��v?���?�O/�$q?���=�?�s?:z�?�٪,-H?Q�?��?7B]?m��?��?J��?d��?��h?X��?9~-$��+c��?��?*�v??>q?=��?�ћ?�@�?J8n?��7=��??��?��{?�Ӎ?�*�-L��?ŗ>ɘ�=� �/^�=R��=E'�,;�>��,��=�q�=.�},"��=.<���+��=.�>�M�=� >Aq>>_�>�X>���=О�=(j>L� /z�>~.:��=-[�=��>�.���=��;׶>P$�=([>���,���=#y>>Z��=u(>��>?U&>m>���=��>JJ-oǉ+�A>&� >� �=�l�=ކ
>�.>��>*A�=bG;�m>U�
>���=.>p�B-�>��?`�S?�΄/ �N?�S?�/G-Z�d?߻�+��Q?��S?�v�,gFH?��>M��+˄R?�}?;]M?��]?X��?+�^?!�u?�2?NH?PZ?5��.��f?^�2.a�R?��N?p6�?��/A7P?�#�=��`?��T?t}?a��+�*?(k?m�b?x<?��s? s?�/�?�c?E2A?�'}?���,(3e,��b?V�^?�rP?N�N?0`?��?<�]?��I?� =\p?l�j?(JM?�v?�i-34�?F�>���>���/�/�>��>'��,>��>�,l|�>��>�h,���>��l=�6C+Tj�>���>��>���>�S?Z��>;�>���>���>�>�;/��>`8.�>���>d:?��_/�\�>���<MB�>6X�>�T�>?��+���>��>p��>���>`4�>�<�>I�
?0z�>�5�>��>I�B-�;�+@�>��>��>.�>��>7��>l9�>���>��<~��>�7�>U��>|��>�~}-���>�I�(:��,6D,覧,��+�� ,3_�)�M&(�,y&��,��'�Gy'F,D��,�J�*��(��,'�+�e�+d�x+�ٛ,8�,J[�)X ,�Ձ,��,��+��':W,y�+��O'�`,I�+��R,��"+{��,S��(���+�E�*O��%+�w*�[�+$��)�,�+��5,v�W+^��+i��*ߙ<,= ,'�&톭+ւH+�+�p�%�9�+��c+D�,o�<'��*�RR,nc�+���=�=OD.�?�=���=R�,+J�=��*4M�=ձ=4w�*�%�=�<<��`+�G�=s[�=a��=���=?�>���=���=���=�J�=��=�.�,�3�=�vc-�3�=Pƭ=8#�=
�r.Ky�=�t;�H�=|ַ=�0�=-ƭ+)��=Z��=�A�=�=a�=_q�=.v�=�5�=�X�=:��=��>,v�j,p��=�ҿ=L��=<Ǻ='��=A��=B�=�*�=�j ;)X�=��=� �=��=�),#-�=��:?��?�)�/km?6?�s1,�u)?V6�+�2?Ӌ?��*�'?*3�=�*,ѓ?T�;?�?��#?��q?I�'?:7?(�?dZ?��'?;O/@�0?^�.�=?��?��=?�i7/��?�I=�)?�s?��4?�|,���><-?�Q(?s�?��5?^�2?�aW?V�(?�a?�8?a!�,�L�)W]*?�N!?+L?�?�)?�Y>?Ns#?X�?���<��+?��+?�=?�(1?��P-�O>?�>H|�=�w�.{0�=�L�=E�,�*�=m��+���=5y�=�?�,Q��=<���+���=���=@��=���=�h">���=dp�=rG�=6��=�g�=�=.G�=L�f-2Y�=%:�=�=C3G.X��=�|9;��=H)�=���=��,��=��=���=iߤ=4��=���=t>���=m��=pr�=�v�,�A+���=m��=���=�b�=�q�=&�=��=���=] ;��=�r�=�\�=g��=�+,]�=�R;?��?Ï{/jf?H-?�F�,�
#?��Z+,�?ɬ?8��++�?v��=��0-%�?�3?2K?�?��f?�#?��0?�I�>Im?�Z!?�I�.��-?�+.bi?!�?��<?ܛ/��?|
V=!7$?B#?T6?J}�+v��>�+?t"?�?�7'?��.?�@O?�e#?��?�)1?&o<-)_�,m�&?7�"?0?��?#&?��6?^]?'K?��<�(?�)(?�?�k,?��9-W9?��H?g(?�/�g!?C�&?�4-3C6?j��,f�'?�%?^Y9,L�?~(�=;�,�$?��C?_&?׍/?��|?��3?*^A?��
?]?�a4?�7/�B7? .F�(?O!$?~�L?�/�?4ES=<�0?��#?ʌF?��+��?�'9?N�1?�^?7�;?`:?�<`?�D/?U?�7E?2��-�*_!6?Ny,?�|(?h$?kx2?�iN?�:/?U�?���<��4?GL6?��"?B<?$�`-�GM?��e?"[<?7/0׆5?ϧ=?�O"-��N?�. -	�:?��>?�D�,=0?؆�=�2,&=?��_?�=?Q�J?��?Q�G?�BV?��?��/?�I?�p�/n~V?\5.q(>???�f?hB/�5?=\|=��P?�6;?��^?��--?��P?��G?#?�hU?�ZW?��~?z[L?��2?�d?�R.�Gq,VP?�tC?D�9?`9?6P?M&e?[�@?�e4?�=mL?|"M?�,<?�aQ?t��-��c?E��=n��==�.�\�=�@�=���,aV�=�$+ղ=/��=�{,
C�=E�;���*֌�=!/�=G�=e��=�Z>qN�=�9�=h�=��=���=��-��=�%-���=���=���=�:.5��=N;��=b��=JE�=0#�+�^�=��=���=f��=[T�=��=CZ�=y�=�Z�=ĭ�=ہ)+��+���=8�=3g�=a�=b��=Z>�=UP�=ň�=;zx�=��=���=b��=-,���=Snf?9?�9�/��4?�
8?L�V-�fL?8F�,��@?��=?��+~N1?�">���,��=?��Z?��F?�)H?c��?�!G?<}[?�� ?�5?)�J?�0
/(~W?��.=?i/<? m?n�B/��1?=p�=|zK?��5?:�b?~S�+�K?9�R?<~K?�#?�JZ?�V?���?åN?'�4?"�e?��-8+�H?��A?n�;?�9<?�R?@�b?��E?��4?c�=��N?�S?|`>?�?P?�ߢ-�6g?e�~,�n*(��*��+�7�)ȹ�+��*̔*��	*���,_��*���,BSV(���'�B�*�Ŵ,�M|*�J�)_8,]E�,IG�)�#,��*&��,Eu�)Sc%*�)��+�4,� 1)\L2+U��+`S�,[ �,���(��t)���,4�+�$+�Y,�5+e�*zQ,���,Ǯ,�w,L$�*M9j*ǭ�)R�,��)=f*�8,�M5+8�[+���+=�+��,�Q+o5,k
*?�,rd,��})���?e�o?��03�o?��s?�_�,&��?#,�o?��r?<Ԋ,�d?,�$>5��,��s?�)�?Zsr?=x?N�?ο�?�B�?|�K?S�b?�3�?_&/� �?tW./�p?��r?t�?�Z�/;Vk?��=;8�?DXs?�<�?�b,�?F??U�?gGV?(��?�F�?�R�?���?��b?��?�^�-��+���?Iss?�Ho?�xk? ̂?Fo�?�x?�']?�R4=���?��?��p?���?��-s�?	�>�-�>)��/���>j�>e�-���>��+<Q�>jR�>�*-Zv�>��j=x�,��>�U�>���>���>��?�#�>;(�>�>���>���>��)/@v�>�8.�Ѽ>Yܾ>@�>�/��>w��<���>��>j��>��:,�B�>�v�>���>Qí>�[�>.m�>��?{T�>G<�>�v�>C�,;R�+n��>���>�>�D�>���>���>f��>��>h�<��>��>r��>8�>�B.-��>�z>1�=DJ�/"�=���=0�-�;�=�;�,":�=|t�=���,��=�i<��+���=�b>E�=G��==->���=���=�:�=B��=0U�=�P�.3h�=2T�-�=7�=�#>�T/W�=T��;5O�=P\�=��>�z�,J�=���=1��=�v�=�0�={�=:>�,�=H�=�>��,��, ��=x��=��=��=MF�=#�	>kT�=,�=���;��=Z�=�i�=q>�T�-�!>&I�>�RG>���.] G>,P><p_,�/^>(Z�,G�E>$LG>���,�:>j��<�A�,�C>�Yn>�MI>W\>G��>��[>\�l>�,>�A>�R>�ak.o]>�Q�-�0I>�B> Ct>��.w�?>�1<�xZ>�'I>��l>��0+v'>{�_>��^>Y�*>7�f>P�h>�ڋ>B�M>�7?>�qn>�B,w�+$ve>��O>�G>�C>�de>�y>AfY>a7;>��;�R>�D^>]�K>\�j>�-��s>>_�,��+f�!,[J.-�6*AfZ,yLT*v�,���,�B�,F,��+Yr�*���*��(,��,��)�y�,s�*��*��,�B,�d,X�*iV�+C�(kF�,�w�,4�+�@�,�4$,S�+�Y�+٥�+x�=+�3+�I6%y],H�L,��f,��')��+�M�+�ʠ(��,�}�*��W,�H�+-M,��,6�;,�}6,Q�+�f�({�*�+3d *�`�+š4+�!,|��,��S,|)+��R,|B@��?x6�0�Q�?7��?HT-�4�?Gˏ,|��?d��?�� -�=�?��>9�:-k��?$��?���?ߨ�?$&@oa�?���?�0�?�?���?��/���?Ĕ/���?3��?z@Ɨ�/gE�?n>\�?���?>?�?�9�,�d�?U�?ZY�?˨�?�?�,�?�@���?��?ջ@�.�3�+G
�?\�?��?vz�?��?\�@��?Bc�?u��=Q�?_��?P��?e�?�ۼ-�@�l?�y;?��0ϱ:?l\A?5W�-g�S?�2H,B@?�X@?-��,��:?�>Aڏ,��??Bh?ߌE?*�H?Fԗ?L?R a?��$?OS9?��U?��/ �W?��g.];A?GYA?��p?	�9/��7?ŉ=)U?��B?�2h?ѡ�+y?�1T?�5P?5�+?o�`?M^?���?�7R?zl8?Εf?5�}-��*uT?]�J?5�@?wC?��Y?�p?��H?i�8?��=��W?�AX?�F?�6b?s��-�o?�d�?�Y|?��/qGw?�Kx?�\-^O�?�z-_�{?b�|?9g*�j?�,,>=��,ʝ}?ڦ�?=U|?t�?'	�?��?ll�?��U?��r?�`�?S��.W��?X�E.� |?�x?/̙?��&/`n?���=��?�iq?���?�&
,��I?ur�?
�?� Z?p-�?Ō?N�?�	�?��o?�A�?�g�-�}�+��?y�?pHy?ʬs?#�?���?Y3�?��j?fKH=h��?�É?pX�?���?�u�-�A�? h�?�lu?G��/ESu?�9v?�_-�ˆ?�g�,�Br?Hoy?���,��f?�K>v&
-�t?�=�?�Pv?y<�?܁�?�<�?��?#vK?�>g?��?�T/�Z�?�v.R�x?��p?})�?O)�/nl?'ϝ=巂?��o?��?�Pb-~*G?	Z�?�σ?�8Y?���?ͣ�?4K�?��?�d?�$�?ʰ.x-�+wv�?��{?8 u?�u?���?�ė?��|?�g?��.=�Ć?���?z�o?��?ͧ�-�>�?�Ph?��3?�/45?�3?��-�?G?*�n+�7?=W7?��o,
�+?�J�=��,�,6?��\?��9?FA?)�?jF?ofR?12?�,?E�B?ئ�.�`Q?"!-.��3?��6?<�a?^�F/?�-?9�y=��K?28?.i\?F��+�P?-M?�'>?vx"?�N?K_O?.�u?o�D?*	+?�Y?���-i�{+�iB?kA>?��2?0;4?��C?f?e'>? �,?�,=�G?1gL?��;?��Q?=�:-��`?��?�o?�W-/��m?�ks?��P-��?Ș�,I�l?-=t?�y�,�+f?��>EHo,X�t?�u�?�)m?�@{?彺?���?k��?�WG?��f?.��?=�A/�Ǉ?��.jk?��m?��?��k/�f?�D�=�E�?�n?��??��+��B?P��?��?�P?3�?Pۊ?R�?��?�4c?�Ӑ?�-�h)�d�?�8y?"�m?.�m?�?b��?�~?�h?n�:=��?�?h�n?�K�?CS�-s�?��?-�u?l$�/�q?Iw?*:�,WX�?E��,�Aq?��o?��5,}�f?�>n�+��w?��?�p?�Ӏ?���?;��?亏?�dJ?]�f?l$�?Wc�.��?ņ.Bq?��s?��?aI6/�Fj?Cߠ= *�?��l?���?a�,inD?�Ŋ?ӄ?3�S?�0�?��?Dh�?C�?�hh?=��?�� -�,�ނ?v�v?@jo?�-o?�[�?��?�<?wi?��2=�7�?��?�v?�6�?�z�-;��?��?B`�?��G0Qß?R�?�7�-��?��-;�?P��?�R%,ى�?��X>s��-�I�?#��?���?B�?+��? ��?g��?@�?E��?G�?���/�ڴ?� �.���?~�?���?8�P/@ݗ?��=�S�?aO�?�B�?�M�,���?�´?T0�?�Վ?e��?L=�?��?�r�?�K�?�ո?U�i.�J*,�ۯ?��?���?]��?K	�?���?�?
�?�@m=��?>0�?�!�?�F�?���-���?�ܟ?a��?e{�/?Do�?���,�I�?M�+�΂?o��?�c�,��?M�4>��.,m~�?�?�A�?]�?!w�?�Ս?p)�?Ќ^?K�~?r�?d�/�%�?�l.t<�?h�?}c�?9:/(�w?��=�	�?-�y?���?���+�jU?��?L��?�Cm?7�?���?Դ?4ڎ?\�|?�̖?��\-yݬ,sS�?R�?s]?�N�?�?��?�7�?�cv?B�?=}��?7��?��?��?��-�I�?=>���=l�$.�^�=�\�=1I�+&f�=�7�*���=2��=qh�,g(�=2�<��p,���=;�=T��=)��=��'>���=9�=S�=4��=Zl�=��;.���=��P-;�=Wx�=�� >�"..���=U�a;�{�=A�=�s�=��*yD�=���=[=�=!Ұ=5��=*��=*>77�=]:�=�� >Ҹ,���*�Z�=O�=��=ӕ�=z��=�S>T#�=�y�=!�;�g�=,��=��=�>�lr,��>�?р^?��k/\?,�]?��-G�v?��P,.�b?@_?��,�'U?U�>*N�,�Kb?M��?�^c?�n?��?�8o?(�? <?:�Y?(�s?2#*/ے�?"z+.�vc?,_?�ى?��_/3�]?m#�=��p?+]?=L�?��,�W3?uA{?�ms?w�C?T��?�|?��?ٔu?��S?�p�?N-�i2)��o?��g?p5`?]'\?4�q?��?��k?��V?��3=fy?�{?��a?�/�?_l�-aY�?#:?�?c�/(�?Jw?0K,�#?'lN,[k?�?���,8�?��=^@�+��?�w/?r�?��?_o?�"?��-?51�>	?�i?���.�$'?)�.n?Z�?>59?*(/�;?^9=8�%?�<?0?���+N�>�)?c�!?oG?+?d�*?�`L?�� ?ӽ
?��5?8��-�1=,%!?A ?�?�o?��?��6?��?ݲ?f��<J�$?�'?��?�T'?���-��7?��?O?70*lw?9Fy?! -�Ɔ?tL�+�	�?�yw?@��,^�l?�c%>���,�6w?pے?{�z?$e�?c��?hT�?>��?��S?�^n?B��?��/G��?�}J.%}?Brz?�ޙ?͢8/l�q?�+�=Qe�?LIr?4X�?7|n,��J?ڶ�?B�?��[?3��?}<�?�?�?�R�?;�h?�o�?��.	�#,�ބ?X �?[w?ٟt?�a�?:��?f�|?7�n??�<=��?q��?�nz?X5�?8�Q-�җ?���?I�?��/L�?�ב?�#-��?���,Ij�?(��?qʜ,���?�C>>��-jV�?d5�?'�?�?���?�؛?Y�?Q�o?B�?�ŗ?��5/�&�?c9�.[�?	e�?��?|/�?s��=�?Gʊ?�C�?���,g�f?�?3@�?�|?�:�?d�?�=�?+'�?�$�?J��?>JU.*P,.�?�y�?6�?P�?��?���?0��?�4�?O@[=$�?��?0��?��?�|.^ϲ?vB?��>��/���>�(?�j�,�4?�w,���>�d ?�,w��>�=#�+3�>��?���>mi?�,I?{�?�?���> u�>�?�ֱ.
?��-�u�>�L�>;�?]�.���>�'=�?
?p��>>�?8�,t{�>W�?�Z?Xe�>��?C�?a�.?(\
?���>c�?�3�,ה�,Sh?�?�T�>k�>C�?�-?8?�G�>�l�<�?vo?�>�*?�b-�Q?=��?�1�?:g'0�N�?�.�?��V-�|�?9:*,�?�?$i�?�+�,FP�?+7>O��,���? :�?�c�?���?��?C�?�7�?��i?�ɇ?���?�o/ib�?�9).��?�J�?�q�?��/$[�?+��==�?��?o��?�,��b?,r�?Xʕ?a�u? ��?{�?���?�n�?��?aЧ?���-Q�*"*�?�v�?Z�?br�?��?y��?貑?���?��Y=�!�?+��?�Ì?�z�?��-�Ϊ?�
>�U�=��/���=C8�=��-�X�=%��+��=TO�=PC ,S��=�#\<b@�,|P�=_Y>��='
�=�{)>/^�=zw>콼=���=��=B_�.<��==!#.�=���=	>r�M/<��=7��;�V�=XA�=�
>��,���=k~�=�-�=�Ⱦ=1<�=��>#�>C��=�L�=� >B�-��@*��=���=�v�=�5�=�U�=�'>���=�N�=h�x;�!�=�,�=X��=�j>��u-�>�+�?�X�?�#0v�?�\�?�S-�T�?I&5,rщ?˃�?}i,��?M#5>��,�d�?��?SW�?�?V��?���?q�??g?�x�?�n�?]v/��?n�.�R�?O,�?���?�|�/P��?Y@�=�o�?*F�?�/�?&N�,�h_?q��?���?�Wu??��?>��?Q�?Ɋ�?PX�?���?�l%.g_*R��?�8�?��?�ދ?��?�?�?
�?��?��N=ZӘ?��?�2�?���?>�-��?���?�B�?7�]/Ҵ�?�s�?�-�t�?;��,�Ї?�?d�w,�y?��0>�yE,l_�?��?\�?�?M�?���?��?td?"��?P�?y�"/5і?�#�-��?K�?�l�?�1#/V�?���=*#�?(��?r$�?�,-�(W?��?)2�?'2i?���?��?���?O��?>y?��?l(-.�)��?���?�M�?���?{��?Bӥ?�?ex�?M:J=wE�?ǔ?��?b�?.�--��?X�?���?>��.**�?��?b-�ގ?W�,?I�?J=�?Q�+,k5}?��0>�ǣ,9�?��?�Z�?J[�?���?�c�?�_�?�^g?�?1v�?1��.�l�?T/K.�ʆ?��?���?Ǳ/��?�K�=8��?�փ?2��?�c�+�*Y?�t�?���?8j?
q�?o�?��?�ӑ?`�z?�[�?��,���,#Ǐ?堇?���?w��?��?�D�?�׌?�^�?"�M=T-�?��?�׆?/��?��u-�y�?qK�?�b�?���/I�x?�k�?�f-Z1�?��+Y�v?��?1n\,sKv?��,>@��,�|�?��?7l�?��?��?���?H��?v�S?�+z?�-�?jS1/ B�?}�-��?B?U�?��"/��}?��=a:�?$�?1��?�x�,h4S?\��?�	�?	�e?w��?�?&�?FЉ?3r?�9�?��-�K�*y�?���?��?��{?��?њ�?���?��q?��E=f��?2�?�w?��?�-fw�?2�?]B�?٫�/�	�?�ŕ?��-���?�Q�,�7�?}��?ǼW-��?w�N>%N�,���?���?�?)�?�?���?�?V^~?���?z��?/:/@��?�iv.��?�k�?Qڹ?5��/Z��?�f�=��?�~�?.��? �*-�ns?I�?���?X��?ZZ�?妥?�?;`�?]\�?�;�?�w�-���,��?z�?'��?>Ȑ?���?Jw�?
'�?�&�?�j=l��?�c�?&�?���?��-*�?��t?t{N?���/4I?BNL?Op -��Y?Oy�,��S?�L?7��,�6B?O�>�o-ǍO?E5s?�8N?tlZ?*Ǜ?�Y?�:h?��*?-N?�]?iM/.df?/	.ǭN?hVM?h�|?ܢ0/KK?p�=��]?P�K?��m?���+]�#?r^b?��]?9�6?�Vg?�Yg?���?g�\?��A?32x?��,�Q�*��a?KSO?qL?��J?�1e?/�|?K�S?A�D?�=6�a?��d?{O?Bq?+K;-O|�?|�7>yT>4�.�>�`>':,�#>�E-��>Z&>�r0,�>���<|�h+ߜ>�0.>��>6h>W<W>ߺ>M+>DT�=�t>Q>*.�,!>'�d-�>>�2>��.`�>���;k >�>�Q,>�^+
��=�">�!>ת�=�� >Y�&>j�F>��>&p	>u/>>m-��(_�!>�>��>��>ڪ>"�*>cp>T�>�ʑ;cX>��!>2E>��*>��,��0>���=ϴ�=3iB/�
�=�=��d,���=�Z�*g��=��=cd�+�6�=B��;�,+��=S�=���=��=[�>:��=b�=FS�=���=*!�=�.t��=~R�-ᬷ=C��=���=][�.�ܲ=�_N;���=��=˷�=+��,=F�=\�=���=��=s��=�;�=�� >��=��=�S�=��-L@�*$��=d�=i�=�ڸ=�4�=b,�=N��=ꃵ=2;З�=zO�=3��=5~�=��6-���=y��?�[�?78�/��?�e�?�YQ-��?qI�,I�?w��?VX6,���?!�4>��,JS�??ވ?�;�?�P�?�?cM�?i?܃?�ڑ?��.�7�?I.�?J&�?���?!+/A�?1>�=�?�?'�?��?��+�_?#�?�F�?y?�N�?ǋ�?68�?b]�?��?أ�?���-�`+���?��?��? �?�*�?��?o��?��?[nK=X��?ZF�?S�?:"�?*��-L�?t��?�v?��/�tr?(�s?V�,)�?�+r�r?݉t?�\,{e?ܸ>��w+p?��?��t?��~?B�?ʳ�?���?�K?��e?Pӂ?�x�.'�?��Q.,�t?XSs?#�?j�w/Q�j?%%�=�@�?��p?�d�?�q<,@�G?��?�\�?tT?�G�?��?~[�?��?Ld?.�?`��-ש�*��?ږ|?��q?H�o?�&�?.ʔ?Vx?b_e?-�1=i��?Br�?hBo?E��?�z�-� �?�Z?�/?|�5/�.?�H0?�-�+C?��+}1?/?��-i%?��=|,�0,?5cR?I�+?�:?A��?��=?\�H?�?�'?��;?�/��C?���-YO1?o�0?Z?YQ%/B\-?�``=��>?��0?-�S?Ir,rw?�GD?�8:?	%?�E?slE?Y�p?Yv;?i�%?�P?�l2-ʧ�)r(B?�08?n2+?ٔ1?AIF?uZ?�m7?�^+? =�D?��B?Җ,?�E?���-��X?f�Q?7�(?T�0)?n/*?y�-e99?��t,O�*?T�/?��#+�O"?��=��-J ,?~�I?�v'?o5?1ρ?�o9?��D??x?9#?Ok9?�r,/=?Ƅ�.��(?�)?�T?�=D/g$?h�m=��1?T/&?��C?�,��?�B?��5?�?3(B?df@?�-i?ƻ9?/�#?9CJ?�H�-�H+C�7?�5/?�1*?&&?��8?�1Q?Z4?��?��=�:?��=?�)?��A?5��-��N?{֚?5�|?ٚ�/Wy?��?�ù,/��?��+�{?���?:T�,2)u?3�)>�9,i�~?���?�-z?�3�?���?���?S��?��W?Aq?gԉ?��&/I,�?��.G�z?a~?ߌ�?ΩH/�|?���=J$�?�? ?�9T,�(P?��?@�?ҋe?���?�N�?d��?�?��s?.w�?��,��,�0�?ے�?�e|?��q?�s�?�
�?_��?Žq?L{9=�0�?3��?o}?%��?'-�?                       @       @                                            0J                    �                                                                                                                                             >�d������}/�:���4
'�ke[#�,;���{"�>��>��nA;��⾾�T��,� KP�5!�+K�> �	�
�Ez��8�:��v�pb+�t��]�F��Uv�=������p1缳?����E�ѪI��wо�?�����w �ٸ"���/���7��M�{tʙ��%	�r�þI���9��9�)��^Z�]t��J�9�����;LT��O�h�þ�n��ƾ        0       1       2       3       4       5       6       7       8       9       10      11      12      13      14      15      16      17                            SNOD  (       �@                             0       �C                             8        G                             @       �                             H        I                             P       (M                                                                                                                                    @       @                                            8N                    �                                                                                                                                             ͋�?���?S�	1d��?Ol�?0�E-���?J.o�?��?�{.��?���>H��.�Z�?F��?��?���?�)#@?��?ȕ�?bײ?���?6��?��K/Y��?a�/���?���?�@є/�B�?%�>d�?���?~#�?��-,ĩ?!(�?VA�?�+�?��?��?�@�*�?h�?4� @��/0��X-���?R�?}��?�L�?��?yh@���?'B�?�7�=01�?(��?�d�?Y �?I��-�6@             (          @               @                                                    HP                     x                                                                                                                             ^I�>�
&q�>��jQ�>2�>��>yܚ"�>��R>��[�2�>=�
?��-�	�qR?:��(b�>2�?�R�>��+(�X��>L��><�>��>�7���	?��?F'�>!����>b���\D�B�,vzD����,��=�1���0�r���<C� ��ХZ�ec'bo���L����� ���N�l�6�H*,}s�H��z�@o̽<-��Ϻ(�]���M��5����h!����<�����|���os���>��Ä"|�NI�� 4=6���1�������W��X�Gs�VS�Z]������j�Bo&�HCF�u���]U�?��tT���k4:����-N������0L�X���L����mv�k�-�4ν�++��_�U�I�J�'������)�D��"�#�����޽X����p	����$�/�$J#���������Vz��7�d䣾8:����~���PE�57���~u�����7���b�DC���k9H���ɨ������W��D����_���,v�f���]��:u�Z'$�"��������d���<�x��rU���$�mׄed�5�g��E���c
�W杄��^��Ӄt����&)�m�Ha�ɰ�xD�+�J!��n0�&Z%͡�=��_�s�mӊr�Χ^�*$�q(+�v�6�f�-�U��0��D� ���y�����G����q� ��0`Ƚ`�&���1����,�2'��4�&�X~��O.����8i̽��DꕽP����T��\%������v����L���)��.��0�z��18��d����Iv��
��r]�Y��a�h6m��P���R������[�Fۃ�I{�͜�O�d��%̓���G�G(Grr�PJǒ-��7��A'���\�fՀ��*��C����MBL1$��X�����l�r�wr��`�P�a�1����2�T/j�T�R��B�A ��!��� �k�t�C���H|r��w`���%��1�37����������־*��1	���й��������?�����+� �䨒���辥�r�_���۾�B��d)���U�=@;"�p��@����?����\��7���Z��V�9m߾͙���r���M�TK�Dnź�?�I��J���槄�� C�g�K��ӊ���1bפ}>�ed�˄*�y�5al�r�/�(	5���F��H_�\U��(�;�+V��!��f#�&$mimK>�xK��ø����v)ă�K����ٽ,���*x. ש� �C�K��P������'/�w7����j�!&�ǽ�< �p�콚G᫇������xV����v�� Ͻ���dK�w������� ѽ~}��F$, ��E+nd��e �̵��[�f�Hx� �l���"��!ֻ��.� 5��mڄ�'�D�����~�)�����:M����ջhd뻂���:��-�s�ie0�i�(��������@��l��B�Ԅ��a o�U+��\n��i��3��k&��Y�Z<�2�,�u��f�X
\�b�e��%�TޱǄ�`auIS���'�����N�d�V��m�dX($Dj�V�t��s��������E�����t7c���6����B��)~��aо�:��:��[¾��)r@���Cɾ�б��������/�������]D������i�,�Ͼ�&¾ga����)2Ş� =�=C�c�p��=��:�=���=�|�=q� ��=HPG=� �P�=0� >���5���H��=W����=���=(��=�r_������=((�=$B�=�C�=Ҋ�pC�=���=@��=��K���=�h�vh��`�����}e����W3���`l|�=��`׾*���i��I	> ����'����c'�G����g������2ؾ{��5'��aU�}�	5�+�!"���S54ʒ��N���:�����y� ���0U��Z�M��'�_x��|�����f�<���j-�$k��*'����S��lf�����Q��$f�|�u�N�(��N������h��"z�����������_�a�p�^��W���ES�]_�2����0�G�2��T���_\���E�����<X��[C������g��v��8���Wߣsjք{�H��vW�(�7P{��c�1a��H���/o]�ܽ�Gs� 6�l����D�!AH� �i@��"�^�@��0풼� q�� �0S^�͙�'[� Z�W�g��]$�Яv��B��MR�&��p��*	��mǼ �5��� �l�p�e��[�m�  �e���#̈́-躾��,�m���㢾�g���d�ǋ�R��3d$�}���̾X�:F�z��	����U��� kɾX�������*V���0����=�����wH�f�̾��¾�ێ�J	��.����	�����H���[pc�(X���ꦽ�K`��Ƴ��{����  h0F{��q���f�;��/ĽGJϩ@��Ȃ���夽]��z� l�������;��잽|��|Žpd�� ̈́�i�p͔�V��<�p�F��"�4��H'��+�(C��@���@��cF��n���W�p�j?l�
,G�����d&��0N�@�6�\c,`�Ft�����Žx<)������Y��AO���ק!� �@�<NZ@C4<GWՄ@�L<@S<@�\<D(`�j<��;�0��ho<�'p<���
 ��O|<I[����W<@�p<@��<��V,��:�;��<��)<@cp<���N�;@<<��o<�f��U<fa�RY�$TJ섄@�[��t�0�w:=��S�\cE�"������b�x6�U������VD�~=>x�*j�
��GR?Խc��"f!g�r8����~�R�Fl��3�V�G���B[��5����H��xd��Y�<܄A�4�нP��B0�v���`��D�߄�X��yU�\lL��Z��̚t�k k�F����5���?����|S_������ю������F���f��]����f���=.���ݬ6���`/��p�7o�D���<��m��pބ�_���9��a��-Y��Z�0+
y�9C����Ԅ�9q�2��z�9ʲ�6����l��w��kt��h����� ����҃,I���󛽈eZ�� 脇��( �����ot������� ���8"����<#̠���U�� ��}�ͩ�u H�m��$��1�LÝ��$������HN��x�����c�1��Z�����`g�3��;����Ӿ�3��n9&�����YD��q{�����M���f���a�>'W��������U㾫Q,�!�eB���W��PVs�DsϾD��t����@����^LZ�ƾ ��<��� =��3 ��<`��<`L�<pSQ@��< �z<5 -`�<��=��� �=D˨��S�< i�<�e=m���� >�<���<p��<�Q�<�+M���< c�<�N�<�Bb�Z�<��X���*}<��k����r0���p<���ׄ*�
�_1�I!���� z�Yb��c�';?��Ed?���W�[��w#�;Y��U!���<{a�Y*�AH�h%�����8�"��ȂQ��d�@�'��?�,���:5�����7:����m�&������W����(��'��Ze�DhJ�[�-������42޽�V9�I�%��)o�P2b��7#�u��/��!����?��{ͻ'�W�᛻3�����j��č�X�����3n�:��Fw仏VT
ڄT�Ի��m��\��[�޻��Ļ5�B�@��#���H���2:�����EX;����ػL瘻��8����Pѽ�*��������ҽ<�񽸬����ƽ�X�2O`X���������2m����?�"&'⽨���Z�Tè�
����ý$�ý�퍽��񽾍�8�����x�˽�=���L��=}F���=    H�=>�="ɛ=�,!�=
B=i{
��=P�=ϓ�u_����=��(���=�o�=(��=��rZ��J��='�=>,�=d�=x� �)�=���=��=��,���=�i>�F�8��>��`��Tj>��>(:>q��r�\>\�=��DN>,۟>nq8��B}���>*��!��o>�!�>�͋>��:�3.���P>$�`>T�>��>p��<>�>0
�> �e>9�]�z>&rY��W���%�v.&jy��29Ɨ31P��R����1�j�b��E2���[�/��x{���+��E΄��tTV���3���,mb�%j���G�L������:9�˘��*
�'��>'�4��F�>��4�>��>C�o>�2��=�>}>����>/H�>�('��C����>��Ψ��>�>�>�P�,n��Z��>(��>��H>}>�>�$"��>/��> !�>��&]�>�':��9�k��T���8���U��A�a�T5�hý1l���K#��у�G/(���u���{���=�2+����e��̥,���>�"�FL1�@��� �P�S��n����6y�,�9�tKn�G�/��İ���о���������m����|��Kox��x�(�z�
����,�����z�-yԾK�Ħ�#�������ƾ��~����5Ι�)�S�z��K�+����־l䟾ʜ�򵯾��=|�U�;=�w0��*=�{;=���<�,���=P=�<����=��G=vV1Pb ��4=���(�=�X=0�1=�]ᩮz 2=x�(= O�<@�)=�{��p�`= jG=�O=x�`�=������� �ܾ��"�(~���`���U��\")Ҽ��GM2�����M��F��]�������뀦�௾\��tIѾ'�O�m�栘�&i��2�`�������S�l �v|�|���`W�ŷ���>�K%><i�pd�=`�>���=y��ܹ�=���=ƒ(��=�\7>Zٺ�� �$>�|B��'>|�0>�.!>F�F���X`r�=���=��=�>��\3>)> e>?E��>�pݼ;� � ���Jc�`�μЬ � ���F����� �)�F����� 2�Wi�k���x&���Y��~��i(������o�j�P��˼�{ż��]��p�^Ї�pS*�@��@�Ѽ���󼰱
���^P�M�{�O ��'� dϼ:xU���������3����h��5"����<����$��� �G�@=,�@(������C�P� ������S����W�`�A�����S���'"�tD���� ?-����`6	��`��1ܽ/����J��B�?P𽴉C�||�����9�'J[�p�`�A�%�,��,/�@(��*�𱽴 �~q��D�?�hY=��P�ϺD���B"�����O�iEJ-#���=�����M�q�b��0���,*8�(�k��\��@�pYX������)���f�luL��{B�8���,��a��}ҽ�#5��لh\g�Ы\�b�!�8l)�0��	f��������.s�$���i��P��)f����C�������sڄ�G
�<�j^��X�`�@����JiJ���0�ӄ��y�,*hJ)�Pf`��U�����S8*PW���N��W�;�����ք�FF�
:��W�����;�7Â%�q����MG��q? ?�Ny��E�QG�̏�H�p�+z/�����zR��PUW�wةm�1����^AS���H�qFT�G>)�ꀁ>d���J>�b>�w >ᛴh.B>�p�=��22>�&�>�<��%� �>e��4N>b��>�ut>YG�_�Q0�3>8�D>v�	>4q_>N. ����>Ҁ�>HRF>!���Z>�Bj�m� ��y�<q�a���U8���G\^�-��d�3���O�z�����&��ٚ�q�'�fs�n6��D�������N��W�6�a�z���e��U {���j㝾ߴi���'΃��Pz->:HY>s	��3*>�cA>B4>�8P|�&>�>�=�X�>�j>On.�{�� �_>Z����->�h>T�N>D�y(�ZIL}>4R$>Է�=�C>��M��Er>|�_>p�.>�j��!;>Lc��'R	�HU"��kP��~�����ȣ��J�<���D�|��h��X)޽0J1�E�}�:2���&���P@��8E+���0�����`kٽ����$�	��ރ�n.��)�O� g������=<�lS�=υ��=H��=�=�m<�7�=�:=��A���=0��=5Y��(�=�x��:�=p]�=Xg�=��	+Pĺ�M�=�ت=��m=��=�����=-�=�M�=�3r(�=]ص�-"M�cr�nᴾ��˾���
���u���(;�����n��Rh �c�j:X�ӈ�X�q��4��WC���ݾl�)#	ㄸ퟾V1���o��Q̾q��� ���i��O�T �þ���jȄʖ�Ds$��z�nD	�������0��羴|��֣��վ�)��\�-��D(�j�'j��� L&��L�H!^-�s&�\־���h��K����3��9*�p� �/��+�(K̽�Q�*���e �ҽ���󜽨 4���@DU�/ ��s��Lc�N[��L҄���^4���Խ���0P���=�� r=��M���AȽ����Dc彴v����e��Hý��-�����¢��#�U���r
��@���_5�) ܺII9�:=�UǺ�>�Rܱ.�~�����q��4���#�*�b�����Ⱥn?޺�ۂ�����/τ�B��,�9�h4^f��8��=������=�L����=�*�=`�]=�^��b�=�=Ùц=�i�= �"�n/���=�(��`�=H��=��=������=`ǐ=�ME=���=G�A���=�Z�=P��=]�<��=.�Ӿ�q���)ΠӾ�뾤N����6��ǾN�Y���dTA������W���V��		�./�)�Sپ�L��]���~���FČ����Ⱦ+ދ�o����L�i�
���ξ2X75�ྐ���P��S�J(��&��9����0g���� /����@0(��fk�p{<�N%� �H����P3� �T�p�/���+�a�x��*��ɼ�I����Y�0HW����))2����t�=IN���=P2{��a�=�=xv=}�P��=��=�Z8Ɗ=`5�=���,���8��=t��g�= -�=(0�=&��*	�@�=X/�=��F=�Ӥ=�����= W�=H��=�E\���=������ 3��@����iƄ���=�x������u䣄��τ@ZZ�� ף<�����C����c ������;�B���'�p��{hqc����k.�z�,M���,��E�=����=��<��ض=Z�=(�=	�%�ϯ=a:=+��x��=`g�=��[�Ǆ���=؉b'|�=���=0�=M,�J�<�=���=�'o=�a�=:�:�8D�=�v�=���=�^tڻ=             (          @               @                                                    Xq                     x                                                                                                                             ��@�X1_T�@��2ug�@��@hg&@�v�1��s@L<�?� 1+O@�EA���2��/�$�@v9o6K,�@ �@���@�\�6�^1|_T@D�v@~��?�/�@�?j0��A�g�@�؁@�|�0��@��_@�Q1���@K��2zz_@�@qC
@���1n�J@
gj?�!�1|,@��@���2��/��@�36��j@y�@~Ħ@�9�6��(0��0@A&M@v�?Pڋ@�3G0�?�@�t�@��W@d��2�́@̟$0lh�.<�0u��-^u0�[0b��/y��.W0Mm�-+N-�A�/5��0
��-�~<,�U�0 4-��0��0���0��!.��-��/S\0�/�2]0��,�+�0L#�0��0Z�,d*Q0[�)@�F�0$щ@�b�2��)@yV@��?�R�1�@�G2?i�1߱@���@��2�\2/ć�@2�16�72@и�@(}@�֤6Ҡ�0�@L�@E�?�QT@s\�0��@�ڕ@��#@l�02E@�fL@s�u0�¥@�#�2'L@ǀ@���?ô�1 29@��V?��1�P@���@=��2�n(/�7�@��]6�lV@��@w=�@}W�6���/zS!@mu;@�/�?f@qE0���@'5�@�=E@���2Ym@Ѱ�,��m+k_+#u)�k+p�i-r�-�N�-w4,;-1,1"*=x�*s�q->x�(2�)-�X-�ɉ,�+V��-�u�-X^,�/*/�-�!-��*-j�
+%,Z-T��+��T,[(�+G�,$B,��,@���0N9�@x��2��,@�Y@6��?��(1�@�q5?���1t�@��@W��1h0N�@Kt'6�W5@��@aɀ@�m�6�;0�e@ހ@�ٔ?�X@��/�Ъ@/x�@n�&@7��0��H@���-~R,Y��,�+ס�+���+�2-p��,=mZ,vN�,�0*��'-�Ӂ,w>�-i�D)���,P�*!O�*DT -�e-���+��s-�2,��`-���+��?-^�(٩,(^�-ņ�+��-4zt,�@�
�0��@�%2��@�jH@���?�`�1�@�&?�0��?#P�@�dU+D�$/G&�@� D6_�&@e��@!�l@v��6U60	��?H�@��?��F@TV�0�&�@�@�@Or@��i2�z8@��4@���0}�@N�-2��4@y d@��?��1 �#@[�=?���16@���@[��1H��/)�@n<x6M�=@>�@5�@���6��(0��@��%@���?�?b@�C0��@ඟ@c�.@d��0F�Q@��l)�Q-���,��-�g_(z�	*�}(�>�,��-_��+sD�,��,���,��D+~�,G:d-�c,��,^#�,s7�)d�,�?�,W-��g*]��-�:O-� d-f"�-/�N,ZN-+f-ּ�*��@0�0p;~@���2nm@glE@]��?�zI1?�@$?)e	1>��?'�@Z1E�0�'�@@�6LQ$@YV�@�zi@R��6g�0��?˙@V��?��C@>��.���@d9�@�@�L�0º5@Ù�;aJ�-��<ۮ�./X�;���;�ki;6E.-�ڪ;�}�:�5-�+�;,29<#ג,��,��"<(_�15��;�"1<�g<��`2>��,2�;' �;Ѳ";���;i�Y+W2:<�9&<��;�N�, ��;E�O+��-t$F-�/�,ա�,bo�,��,�+?b3+���+�c�-���+Պ-d��* p�(y��+� >*A�m,��-_T<,�,�Q*��,���*$m�-�3-�-��!,8e+�d�+��Y+x��,-�H@�0$Ϣ@�3�mH@��|@A	�?+�1��5@oR?�z�1�X@>L�@�^�2���/��@�Bm6ƂR@��@ˇ�@ǿ�6�;0S@h�7@���?�z@~ӥ0o[�@"�@�A@2p2��h@]�]@���0���@=xO2�W]@���@A	@hs�1n�H@�i?�z�0�*@@��@]�2-x�/�@�aO6{|h@�>�@3�@"�66�0�.@�8K@��?Ou�@�M�/���@�c�@��U@��V2���@W�l@�nK1�ʿ@s��2�Cl@�@�b@�_1�VV@�x?,�176@ W�@�[�1V 0���@H�B62+x@�B�@l*�@3�6�&�/��:@-�X@C�?ȓ@�P�0R��@9��@sLd@�k2�3�@^T@���0��@W��2)�S@���@�"@3�;1�@@��^?,�1f%#@J�@\^�2]�0�ɶ@��]6tc^@_;�@��@�2�6lUO0�Q'@�hB@��?^s�@�k�0]h�@��@!�L@l��2F�u@sN3@Z��/;~�@x�f1�3@Xb@T��?y-(0l"@�;?�h�0��	@FP�@1�<2.o.i��@v��5�<@N��@7��@�*�5��d/�u@�d$@lH�?3!`@a�.
C�@�5�@)-@J`�1�P@�G.@R��0�z�@0��2�.@�[@�O�?��1��@�]6?��s2�@qy�@���2��.mm�@H�O6��6@[ �@�@a�6�e�0�v	@��@rϕ?�Y@]ܔ0{e�@�ؙ@�)(@x�x2j;J@ߨE@SK|0+i�@�2GmE@\"y@^H�?_Md1�3@7O?�M1
@�f�@Zn29}/��@��50_O@��@zS�@P�*6\��0��@ 95@�?0w@_�$0�q�@Np�@h�>@��/zRe@;@���0�˗@���2$�:@�k@�?�I�1�d)@W�C?�X1�@-��@U�1�x�/�g�@*�U6�3D@a��@�j�@�6ӑ*0��@rs+@ʠ?`�i@ʞe0a��@��@�p4@-�0��X@kcL@�z�0�Υ@��z2�#L@�Ȁ@��?�E�1r$9@�|V?�"0m=@N��@zN�1���/�I�@kPc6kV@�'�@CI�@|�6���0?F!@Jh;@���?�r@S]_0y��@�I�@�6E@�v2m@�H@H#�0.�@;�2�zH@�}@?�?�|#1��5@ggR?P��/ed@qa�@R��2 �/�+�@�gV6��R@�ɼ@/��@ƪ�6��0�Z@�8@���?��z@;�f0s�@g�@��A@��2��h@�].�&�+LU�.��+�U.��.�\�-�04-ih�.�l�+<$E*�o.L�'/�he-�a�-q/�&z+z��.lx/���.��F,z.�*4I.;�C.�O�-�ѳ.��-��/�/"QX.��3&��.�.@�q�0�O�@%�2��-@Ms[@��?um�1*�@�6?*�|2��@�H�@�2'�//A�@ҥ-6p�6@�ң@YɁ@���65\-0�J	@c�@ ��?��Y@Ե/�3�@���@*�'@�8�.�I@R�/�y7-�3~/��7+�g�.f5/�7`.���-3��.]p,�8n-�	�."%�/!�,+�Z,���/��+)/p�/��/��,f��+��.W��.ś�-�M/�wl-�z�/#��/ޤ�.��-!�@/�$@��0��@e�e2�#@ԸN@��?s�61Ģ@�`,?���/^|�?�-�@�k�2�Gf/�r�@+l6�,@.�@�kt@�@t6��0�w@�m@�]�?P�L@��/��@襐@!J@��22�H>@��_@b˫0�u�@
k�2Q�_@���@y
@�+1}�J@d{k?�2>@,@���@�s�2z�0=��@� @6]�j@OA�@K��@}0�6�)�0��0@^?M@���?�͋@��0��@�G�@6�W@F:�0�ʁ@�"�@�*�0ظ�@=[�1���@(@�@83"@+�1��m@?as�1�I@%� A��2\s�/�*�@�V	6���@���@�a�@�ه6�Gf0��N@�|p@���?��@
�-
�A�L�@}@T�229�@�w�0�#,Y01�k�,ԩ0%8�0]I!0!M(�p�0%F5.j�S)`.h0*0f1X��,D�k,tB1���(D�0�+[1�) 1�Ɔ+9�,		o0,�0㈌/� �0���,o�f1��C1�I�0(ҁ)���0[�[@$M�0C�@�2,Z[@\�@o�@)��1��F@})g?��1�)@��@0��2߾0�G�@1F6�`f@?P�@���@%�6S\�0�]-@kI@=o�?�0�@5p�/ ��@��@�S@�Xx2+�~@�8B;��-�֝;�}�.��A;Pu;
��:��,��/;LUJ:��-^?;�Z�;Z�'-4�+ӧ;�wA2�K;e�;Y�;��2�%�-�;�2;���:��r;Ng�*�a�;ݤ�;�c;;�SW-*{a;��/@���0e�@��2�K/@Q5]@{�?��1%�@q)8?T�.2�@R��@h��2���/'e�@�P6�!8@��@ǂ@�C�6�A�0~
@h� @��?M][@F�/�v�@eԚ@�Z)@�0}2|�K@�2@�h 1��u@���2M@k�>@ĺ?L "18�@�%?!�/І�?Kɔ@]��2�a�/���@�B6Ѣ@UL�@�xa@iT�6�*�/���?B�
@j�?F=@db0���@�{�@e�@�)m2/r/@�K@�+M0�w�@��c2,�K@%}�@U��?mh�0��8@��U?�4�0��@���@��1��/��@��5�U@�ǿ@��@QS6 �+0O� @��:@�U�?�~@1�0Ù�@%�@e�D@_.22�l@� -]u-��-�Ù*UY-Ό�+~��+��)�~-4+�+dA-�3I)�Ns+~)D*u�-�ݮ,��C+oZ-mF-�Е+{�,�y�+�p�*$,0>�,��,�H�,�X#-��-*�i-щ+�++��R@��1��@_�2u�R@Zф@AB@�x2��>@B�\?4��1"@�=�@�/�2v��/�Ե@��Y6�]@k6�@��@G��6���0�D&@�=A@�Y�?ɹ�@�\0�\�@*��@[K@�Nq2�t@5+@�x�0��@@��2��*@\�W@��?��1��@�n2?'�*2�t@�m�@x�1�n�/ϼ�@�D<6�u3@��@.(@Z۰6U�*0V�@��@��?�U@=Μ0T�@_�@2�$@,"W2�|F@��1@=�0zo�@�܇2�1@qS`@J��?��1�3!@�n:?%˕0��@�	�@C��2��/%��@�76'�:@Qh�@���@���6J��/Nb@-#@��?�y^@��Y0\��@��@�+@�0�zN@��@F�1��|@y�2m}@�6D@�t�?d�1�@z>#?��1���?��@��2R�/IP�@��H6T#@Bh�@�
h@X��6���1a��?b�@W��?��B@�I�/H�@0[�@:@�2��4@�hV@s�1�@|��2�%V@��@M�@�zg1�?B@�Na?��80��$@0��@ᛢ2��/O߸@l#$6/�`@���@���@$�~6�)06)@P�D@}��?o��@���/H��@��@U�N@��-2<�x@�fX@��1/{�@� �2<#X@�T�@��@�e�1uD@R�c?���1s�&@,��@��2�y/���@&<6�c@GW�@�,�@���6���0a�*@�pF@և�?�2�@���0\��@�˾@:�P@�Y2x {@�M@)�W/��}@]f[1�@�E@&5�?R�0S�@��#?T��/�t�?H��@fIJ2�].ۆ@8��5P�#@C �@��h@w"6|�0��?�O@�~�?daC@g,/r��@��@��@uK�.�U5@��'@C׻0
W�@ �2��'@z�S@���?��K1c&@��/?�+<1~,@�<�@�e	1⇮/��@7�,6�80@�	�@�mz@��6�0�}@S @�j�?_�Q@f��0� �@kA�@J"@	 �0��B@�*@+�1��@7-�2w�)@�JV@�7�?7�1*@�X2?S1��@v+�@
t�2�w,/䭒@��I6�`2@N�@$d}@{(�6��0�'@"�@�X�?B�T@&��/��@�@j$@9�2�@E@xL@/9�0S�@�{�2�9L@ڀ@���?H1`29@�1V?�11�D@��@
��2���/�n�@�+%65�V@�R�@Ke�@���6�w0�K!@�y;@��?��@�[�/�,�@�o�@�GE@��e29m@�E)-�~4-;��-or-��
,U�-h��*<�-��-���+���,܈�,���.�ɤ-2)**ڎ�.��,!:e-�[�.�fe.�].Wz -���+�-7N,�n�-Y�+ߪ4.ŏ-��-�W�)o��-B��*=�)�]�-J<*���,�"�,�Cy-�m2*5��*T�S(�ƍ,I�*�e�*��%=�,��3-�l$-��)��M-�+�У,�w-e�,�K,OR�,��x)u�<*!Nk*��);m- 	�+QT�)��\@|*�0��@0�2љ\@-�@�@=F�1�"H@��h?��Z1�*@���@�<n1��.�K�@�LR6,�g@If�@�k�@\�6@�0gh.@�J@⫾?��@ڊ�0��@���@�(U@g�0S�@*E@���0��@�L1*�D@Cax@X��?��h1�2@кN?�UF1��@���@5б2��/���@sh+6A�N@P�@�ڒ@�-�6kK609@��4@E��?Qv@d�x0���@�ܭ@I(>@�h2,�d@�sp@�m�0y��@?��25&p@�z�@��@u�O1	�Y@4�|?�x1�9@3-�@Sl�1Wq�/�B�@ <`6�;|@���@��@p�6mhj1��=@��\@TK�?�2�@\�/Cp�@ ��@�h@���0�q�@��`@�)�0�_�@�$�2/�`@���@�
@o��1*�K@-l?��1q-@:��@��2�O�/l��@�wG6��k@W�@で@�'�6��R/p1@�-N@���?
~�@'��0o$�@:L�@e�X@�Iv2�h�@�qb@�l1Z��@Ҥ21%b@O��@�@�1t%M@1ln?Ѵ31�G.@�T�@���0=��/=�@�63m@��@"��@"�6��40�2@�O@cU�?�n�@$y0��@���@��Z@��A2�O�@��N@��1���@x��2םN@�N�@� @X��1 m;@:�Y?%~0�=@+$�@w֘2i�/-H�@�C�5�Y@�M�@��@�vj6�)�/�Q#@й=@E}�?F:�@�U0�;�@�P�@¢G@u5-2��o@��]@��1��@�i�2W�]@���@.	@5gW1�H@�i?�5:0v�*@���@�A�2�h/E�@�nJ6o�h@)z�@�;�@���6�e�0�
/@dK@��?͘�@�h�0\#�@;��@�V@Ϋv2'��@O�Q@�(�0���@��o2:XQ@��@�@��
1��=@�@\?�N2�I!@��@s��2䶚/�@1�#6t�[@���@ !�@m~�6X��/�j%@I5@@G��?$��@�~0H�@�Ը@�?J@nth2�#s@�5	;ۈ
.7_;��-�	;.!-;�@�:,�F.χ�:r�:U��,���:�I�; -R8n+�8m;j��/f�;%a�;L�L;���1�?,�C�:��:�%k:}�+;V(,+��;��r;�_;�в,,A;��?@rJ�0=��@��2_t?@�q@���?yS�1��-@I�H?���1�m@���@�=1_&�/�f�@OmN6;I@^M�@�ގ@cI�6K�\0�6@��/@��?��o@���/ǈ�@�)�@e�8@Qjb2e^@�Wg@A�0j��@��2�g@@��@E@�sf1ԔQ@7Rs?���1n	2@�8�@L�2��/�g�@��n6�r@�X�@zH�@�K�6��`/�6@r%T@t�?���@|0�s�@���@<_@��a2�(�@�^@	�08�@���2g�]@���@?F	@ �1s0I@��h?��r0��*@�c�@i�1���/���@TB6��h@ ��@X��@��6��0k:/@�K@!"�?*̊@�0Y��@5��@�NV@a2f2Ԁ@&�@@��0�q�@���29�@@6s@���?��1��.@x�J?��1_y@��@�:�2�ы/vP�@:6AbJ@H�@I��@�<�6ܺ�0�J@q�0@�T�?'q@�Y0w��@{�@�+:@'H2�_@L�-_6c+Jx.I�)��H-a��-��-�y�,@`w-�;�-�kf-z�->G[.;��*���*���-���+0�.��.�G�-�ب+˗F,�@-Y7-&�-��-qt)�	.+��-�.n�B(3م-��!@�m�0Uo�@�72#�!@� L@��?��2��@=�)?D�0E�?K�@N*�2��/t@��96��)@Y�@�nq@�D�6�ײ0�x�?Wv@�@�?@uJ@�=�/T%�@P�@�=@�H2��;@                                                                            h�     �               �                                                                                                                                             �r���1��B��L��i瘽a�W�V%����)���o��%���X���C��r�����7#���򥽺�M�y�r�L�[�4�z���>3����=������n���                                                                            ��     �               �                                                                                                                                             �uz<�Y�0n �<~�/�!z<���<V<#-�0�b<��;�6�.��@<���<�0�/[�-*��<���1�Z�<�1�<�t�<KT&2%:	0˻E<��e<A�;�l�<M�-~5�<ԯ�<^�q< �p.�;�<             (                                                                             ��     �               x                                                                                                                             �1q�u��Ȗb�.��HId��S���P�o �|�`��V	�z��4n���g�F#������|�l\�p�W�Xm��-��d�������c�(Հ��9��,m� {��9o��sZ���a�<��(:~�SNOD  h       X�                             p       �                             x       x�                             �       P�                             �       ��                             �       ��                                    �                                     �+                                          (                                                                             `�     �               x                                                                                                                             NR+E�7#1*E` �1:E�#EZfEi0�N.E��WDr|.>�(E�n;E�!.K�/`DE	��69�
E�19E"�RE2a8g�	0��Eږ7EC�D�.Eit�.h�&E� E;�<E�bb-;?E                                                                          �                    �                                                                                                                                             $�˽                                                                          �                    �                                                                                                                                             n�=PK        ! +�M^?   ?              �    metadata.jsonPK        ! t-xү  �             �j   config.jsonPK      (p&Z�n�� �            �B  model.weights.h5PK      �   x�   �       �J@� N��b��R�.