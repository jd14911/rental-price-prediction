���     �sklearn.ensemble._forest��RandomForestClassifier���)��}�(�	estimator��sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��gini��splitter��best��	max_depth�N�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        �monotonic_cst�N�_sklearn_version��1.5.2�ub�n_estimators�K�estimator_params�(hhhhhhhhhhht��	bootstrap���	oob_score���n_jobs�NhK �verbose�K �
warm_start��hN�max_samples�NhhhNhKhKhG        h�sqrt�hNhG        hNhG        �feature_names_in_��numpy._core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h*�dtype����O8�����R�(K�|�NNNJ����J����K?t�b�]�(�Age��	RestingBP��Cholesterol��	FastingBS��
RestingECG��MaxHR��Oldpeak�et�b�n_features_in_�K�
_n_samples�M��
n_outputs_�K�classes_�h)h,K ��h.��R�(KK��h3�i8�����R�(K�<�NNNJ����J����K t�b�C               �t�b�
n_classes_�K�_n_samples_bootstrap�M��
estimator_�h	�estimators_�]�(h)��}�(hhhhhNhKhKhG        hh%hNhJ�
hG        hNhG        hNhBKhDKhEh)h,K ��h.��R�(KK��h3�f8�����R�(KhMNNNJ����J����K t�b�C              �?�t�bhQh'�scalar���hLC       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���Kh)h,K ��h.��R�(KK��hL�C       �t�bK��R�}�(hK�
node_count�M=�nodes�h)h,K ��h.��R�(KM=��h3�V64�����R�(Kh7N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples��missing_go_to_left�t�}�(h~hLK ��hhLK��h�hLK��h�h^K��h�h^K ��h�hLK(��h�h^K0��h�h3�u1�����R�(Kh7NNNJ����J����K t�bK8��uK@KKt�b�B@O         �                    �L@j8je3�?�           ��@              �                    �?�.�� ��?-           �}@              t                 ����?�>ub�Z�?�            �x@                               ����`מ���?�             o@        ������������������������       �                      @               Q                    @I@���t�E�?�            �n@              H                    �H@���mC�?h            @e@              ;                    @G@������?`            �c@       	                          a@�%~^��?I            �]@        
                           �?�û��|�?             7@                                 �l@�z�G��?             4@                                  �]@ףp=
�?             $@                                   F@z�G�z�?             @        ������������������������       �                      @                                  h@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @                                   �A@      �?             $@        ������������������������       �                     @                                  �a@����X�?             @                                  \@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @               $                   �[@�q�Q�?;             X@                                  �Z@�G�z��?             4@        ������������������������       �                     @               #                   o@�	j*D�?
             *@                                �����X�<ݚ�?             "@        ������������������������       �                      @        !       "                   �j@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        %       &                   �c@�?�'�@�?.             S@        ������������������������       �                      @        '       2                   �a@������?,            �R@       (       /                    @E@      �?&             P@       )       *                   hq@`�q�0ܴ?            �G@       ������������������������       �                     =@        +       .                    @C@�����H�?	             2@        ,       -                    �A@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     .@        0       1                   Pq@�t����?
             1@       ������������������������       �        	             .@        ������������������������       �                      @        3       6                   @b@���Q��?             $@        4       5                     F@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        7       :                    �?z�G�z�?             @       8       9                   f@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        <       G                    `@8�Z$���?            �C@        =       F                   �_@      �?
             0@       >       C                    @H@r�q��?	             (@       ?       @                   �p@ףp=
�?             $@       ������������������������       �                      @        A       B                   �^@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        D       E                    m@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     7@        I       J                    P@�q�q�?             (@        ������������������������       �                     @        K       P                   Pc@����X�?             @       L       M                   0a@      �?             @        ������������������������       �                     �?        N       O                    m@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        R       S                   �Z@z���=��?4            @S@        ������������������������       �                      @        T       s                    �?���?2            �R@       U       `                    �J@d�;lr�?*            �O@        V       _                 ����? 	��p�?             =@       W       ^                   �^@�8��8��?             8@        X       [                    @J@      �?              @        Y       Z                   �i@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        \       ]                   `^@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        	             0@        ������������������������       �                     @        a       l                   �b@�������?             A@       b       c                   �^@��.k���?             1@        ������������������������       �                     @        d       k                   �r@�n_Y�K�?             *@       e       f                   �\@���!pc�?             &@        ������������������������       �                      @        g       h                 ����?�����H�?             "@       ������������������������       �                     @        i       j                   �`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        m       r                    @K@�IєX�?
             1@        n       q                    �?z�G�z�?             @        o       p                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     (@        ������������������������       �                     (@        u       �                   �b@�ň?�S�?b             b@       v       �                   (s@
�cՔ��?R            @^@       w       �                   �k@Ȩ�I��?G            �Z@        x       �                   �g@H(���o�?#            �J@       y       �                    a@     ��?             @@       z       {                    �?�r����?             >@        ������������������������       �                     @        |       �                    _@r�q��?             8@       }       �                   @g@�<ݚ�?             2@       ~                           D@�	j*D�?	             *@        ������������������������       �                      @        �       �                   �`@���|���?             &@        ������������������������       �                     @        �       �                 033@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �       �                    �?�ՙ/�?             5@        �       �                    \@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   @b@�t����?             1@        �       �                 ����?      �?              @        �       �                    �K@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     "@        �       �                   pb@�iʫ{�?$            �J@       �       �                    �?8��8���?              H@        �       �                   �a@      �?              @       ������������������������       �                     @        ������������������������       �                     @        �       �                    @I@ףp=
�?             D@        �       �                   �m@������?             1@        ������������������������       �                     @        �       �                   @_@���Q��?             $@       �       �                    �D@      �?              @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     7@        �       �                   �m@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    @��S���?             .@       �       �                    �?և���X�?
             ,@        �       �                    �J@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �t@���|���?             &@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    `@ �q�q�?             8@       ������������������������       �                     2@        �       �                   �h@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �O@�0���?.            �T@        ������������������������       �                     =@        �       �                   �`@���3L�?             K@        �       �                 ����?��2(&�?             6@       �       �                    @J@      �?             (@        �       �                   �[@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     $@        �       �                   pe@      �?             @@       �       �                    r@��
ц��?             :@       �       �                    �H@�����?             3@        ������������������������       �                     @        �       �                   �a@@4և���?             ,@        ������������������������       �                     @        �       �                   ``@؇���X�?             @       �       �                 ����?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                   �r@؇���X�?             @        ������������������������       �                     @        �       �                   �s@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �                       pff�?�6��+�?�            p@        �       �                   `]@      �?9            �S@        �       �                    a@ףp=
�?             $@       ������������������������       �                     @        �       �                    [@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    ^@�ʻ����?3             Q@        �       �                   �e@z�G�z�?             9@       �       �                   pj@r�q��?             8@       �       �                   �^@��S�ۿ?
             .@        �       �                    п�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     (@        �       �                    @O@�q�q�?             "@       �       �                   �m@      �?             @        ������������������������       �                      @        �       �                    �?      �?             @        ������������������������       �                      @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                   ``@>��C��?             �E@        �       �                    �R@ҳ�wY;�?             1@       �       �                    �O@     ��?             0@       �       �                    _@�q�q�?	             (@        �       �                   �`@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   d@և���X�?             @       �       �                    b@���Q��?             @       �       �                    �M@�q�q�?             @       �       �                   �i@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �                          �?8�Z$���?             :@       �                          @P@      �?             8@       �                         �q@r�q��?             2@       �                           �M@      �?             0@       �       �                   @f@�����H�?             "@        �       �                   �e@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @                                pb@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?              *                   `P@8�e����?k            `f@                                @N@��˥W1�?O            `a@        	      
                  �S@�? Da�?#            �O@        ������������������������       �                      @                                 �?\#r��?"            �N@        ������������������������       �                     7@                                �b@�S����?             C@                               �^@     ��?             @@                                `]@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?                              ����? 	��p�?             =@       ������������������������       �        	             2@                                �`@"pc�
�?             &@        ������������������������       �                     @                                �a@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @                                 @M@      �?             @        ������������������������       �                     @        ������������������������       �                     @                                �`@�}�+r��?,             S@       ������������������������       �                    �G@              %                `ff�?\-��p�?             =@                                 b@�z�G��?             $@        ������������������������       �                      @        !      $                  �m@      �?              @        "      #                   b@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        &      '                   �?�}�+r��?	             3@       ������������������������       �                     .@        (      )                  �a@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        +      :                  �b@      �?             D@       ,      -                ����?@�0�!��?             A@        ������������������������       �                     &@        .      7                  �l@��+7��?             7@       /      0                  pb@�q�q�?
             .@        ������������������������       �                      @        1      6                   �Q@����X�?             @       2      5                    Q@���Q��?             @       3      4                033@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        8      9                  `c@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ;      <                  �c@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        �t�b�values�h)h,K ��h.��R�(KM=KK��h^�B�  ���Y��?t�S��?�R�-'��?�Zä���?0�.,F�?��o��s�?��)�?R0���[�?              �?����4[�?3��,��?WWWWWW�?QQQQQQ�?4����?1���M��?�D �D �?Rv�Qv��?��,d!�?8��Moz�?333333�?ffffff�?�������?�������?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?      �?              �?�m۶m��?�$I�$I�?      �?      �?      �?                      �?      �?              �?        �������?UUUUUU�?�������?�������?      �?        ;�;��?vb'vb'�?�q�q�?r�q��?      �?        �$I�$I�?�m۶m��?              �?      �?                      �?������?y�5���?              �?��g�`��?к����?      �?      �?��F}g��?W�+�ɥ?      �?        �q�q�?�q�q�?UUUUUU�?UUUUUU�?      �?                      �?      �?        <<<<<<�?�?      �?                      �?333333�?�������?�������?333333�?      �?                      �?�������?�������?      �?      �?      �?                      �?      �?        ;�;��?;�;��?      �?      �?�������?UUUUUU�?�������?�������?      �?              �?      �?      �?                      �?      �?      �?      �?                      �?              �?      �?        �������?�������?              �?�m۶m��?�$I�$I�?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?        �cj`��?
qV~B��?              �?O贁N�?ƒ_,���?��i��i�?�eY�eY�?������?�{a���?UUUUUU�?UUUUUU�?      �?      �?      �?      �?              �?      �?        �������?UUUUUU�?              �?      �?              �?              �?        �������?�������?�������?�?      �?        ى�؉��?;�;��?t�E]t�?F]t�E�?      �?        �q�q�?�q�q�?              �?      �?      �?              �?      �?              �?        �?�?�������?�������?UUUUUU�?UUUUUU�?              �?      �?              �?              �?              �?        �K��T�?Z}����?"pc�
�?�GN�z�?�	�[���?+�R��?e�Cj���?M0��>��?      �?      �?�?�������?              �?UUUUUU�?�������?�q�q�?9��8���?;�;��?vb'vb'�?              �?F]t�E�?]t�E]�?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?      �?        �<��<��?�a�a�?      �?      �?      �?                      �?�������?�������?      �?      �?      �?      �?              �?      �?                      �?      �?        �琚`��?
�[���?�������?UUUUUU�?      �?      �?              �?      �?        �������?�������?�?xxxxxx�?              �?�������?333333�?      �?      �?              �?      �?              �?                      �?�������?333333�?      �?                      �?�?�������?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?      �?                      �?]t�E]�?F]t�E�?      �?                      �?              �?UUUUUU�?�������?              �?UUUUUU�?�������?      �?                      �?"�%��?o4u~�!�?              �?&���^B�?�%���^�?t�E]t�?��.���?      �?      �?      �?      �?              �?      �?                      �?              �?      �?      �?�;�;�?�؉�؉�?Q^Cy��?^Cy�5�?              �?n۶m۶�?�$I�$I�?      �?        ۶m۶m�?�$I�$I�?      �?      �?              �?      �?              �?        �$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        �a�a�a�?�g�g�g�?      �?      �?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?�������?<<<<<<�?�������?�������?UUUUUU�?�������?�?�������?UUUUUU�?UUUUUU�?      �?                      �?              �?UUUUUU�?UUUUUU�?      �?      �?      �?              �?      �?              �?      �?      �?              �?      �?                      �?      �?        $�;��?qG�w��?�������?�������?      �?      �?�������?�������?�������?�������?              �?      �?        ۶m۶m�?�$I�$I�?333333�?�������?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?              �?      �?                      �?      �?                      �?;�;��?;�;��?      �?      �?�������?UUUUUU�?      �?      �?�q�q�?�q�q�?      �?      �?      �?                      �?      �?              �?                      �?      �?              �?      �?      �?                      �?�l|3�v�?jr�y)�?'!����?ۻ��<�?AA�?�������?      �?        XG��).�?��:��?              �?^Cy�5�?(������?      �?      �?UUUUUU�?UUUUUU�?              �?      �?        �{a���?������?              �?F]t�E�?/�袋.�?              �?�������?333333�?      �?                      �?      �?      �?              �?      �?        (�����?�5��P�?              �?�{a���?a����?333333�?ffffff�?      �?              �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?(�����?�5��P�?              �?      �?      �?      �?                      �?      �?      �?�������?ZZZZZZ�?              �?Y�B��?zӛ����?UUUUUU�?UUUUUU�?              �?�m۶m��?�$I�$I�?333333�?�������?      �?      �?              �?      �?                      �?      �?              �?      �?              �?      �?        UUUUUU�?UUUUUU�?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ/��hG        hNhG        hNhBKhDKhEh)h,K ��h.��R�(KK��h^�C              �?�t�bhQhchLC       ���R�hgKhhhkKh)h,K ��h.��R�(KK��hL�C       �t�bK��R�}�(hKhuMhvh)h,K ��h.��R�(KM��h}�B@G         �                    �?4�5����?�           ��@              #                   �^@n��c���?h           ��@                                hff�?�c�Α�?*             M@                                  @E@��
ц��?             :@                                 �Z@� �	��?             9@        ������������������������       �                     @                                ����?D�n�3�?             3@              	                    �?�q�q�?             (@        ������������������������       �                     �?        
                          �]@���|���?
             &@                                    J@���Q��?             @        ������������������������       �                      @                                   ]@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?                                �����r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?                                   @M@      �?             @@                                 �U@���7�?             6@                                   D@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     3@                                   �M@�z�G��?             $@                                   _@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @               "                   0`@؇���X�?             @                !                   @L@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        $       u                   �`@�������?>           �@        %       2                    �?����X�?t            �e@        &       -                    �J@R���Q�?             D@        '       (                    ]@���Q��?             @        ������������������������       �                      @        )       *                   `]@�q�q�?             @        ������������������������       �                     �?        +       ,                   �i@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        .       /                    �P@�#-���?            �A@       ������������������������       �                     >@        0       1                   xr@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        3       4                   �f@�7�?^            �`@        ������������������������       �        
             ,@        5       <                   �j@���|���?T            @^@        6       ;                 ����?�+e�X�?             9@       7       8                    �?P���Q�?             4@       ������������������������       �        
             1@        9       :                   Ph@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        =       `                   ``@r�q��?E             X@        >       E                   �n@�LQ�1	�?             G@        ?       D                    �?z�G�z�?             4@        @       C                    �?�q�q�?             @        A       B                   �l@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     ,@        F       G                    ]@��
ц��?             :@        ������������������������       �                     @        H       [                   @]@և���X�?             5@       I       J                    �I@և���X�?
             ,@        ������������������������       �                      @        K       Z                 033@�q�q�?	             (@       L       S                 433�?���!pc�?             &@        M       R                    �?      �?             @       N       Q                 ����?�q�q�?             @       O       P                    �J@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        T       U                   @_@؇���X�?             @        ������������������������       �                      @        V       W                    @K@z�G�z�?             @        ������������������������       �                     @        X       Y                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        \       _                   @_@؇���X�?             @        ]       ^                   8q@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        a       d                   `Z@j�q����?&             I@        b       c                    �?�X�<ݺ?
             2@        ������������������������       �                     �?        ������������������������       �        	             1@        e       j                    �H@      �?             @@        f       i                    @F@      �?              @        g       h                   @e@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        k       p                    �O@�8��8��?             8@       l       o                    �?�}�+r��?             3@        m       n                     L@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     0@        q       r                   @\@z�G�z�?             @       ������������������������       �                     @        s       t                    �P@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        v       �                    @L@������?�            0u@       w       �                   �g@P�<��?�            @o@       x       �                    @��;��j�?�            �n@       y       �                    ]@K�(i�?�            @m@        z                          `i@֭��F?�?            �G@        {       ~                 @33�?      �?              @       |       }                   @f@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?�	j*D�?            �C@       �       �                   �l@���Q��?             >@        ������������������������       �                     &@        �       �                    �I@p�ݯ��?             3@       �       �                    �?z�G�z�?
             .@       �       �                   �o@z�G�z�?             $@        �       �                   �[@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    @A@z�G�z�?             @        ������������������������       �                      @        �       �                   �q@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        �       �                    @J@Ԧ\�s�?n            `g@       �       �                    �?�"ZN��?V            �b@       �       �                    �G@����l��?N             a@       �       �                    @D@p��@���?1            @U@        �       �                    `@@�0�!��?             A@        �       �                   `p@X�Cc�?
             ,@        ������������������������       �                     @        �       �                   �e@      �?              @       ������������������������       �                     @        ������������������������       �                     @        �       �                   pf@P���Q�?             4@       ������������������������       �        	             .@        �       �                   @b@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                    �I@        �       �                   �^@      �?             J@        �       �                 ����?ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        �       �                    �?����X�?             E@        ������������������������       �                      @        �       �                   �q@ҳ�wY;�?             A@       �       �                 ����?     ��?             @@       �       �                    `@���N8�?             5@        �       �                    �I@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        
             3@        �       �                    b@"pc�
�?             &@        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     &@        �       �                 033�? ���J��?            �C@       ������������������������       �                     B@        �       �                    �?�q�q�?             @        ������������������������       �                     �?        �       �                   �o@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   g@�8��8��?             (@       ������������������������       �                     &@        ������������������������       �                     �?        �       �                    �D@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �M@���R��?6            @V@        �       �                   �h@r֛w���?             ?@        �       �                   �e@z�G�z�?             @        ������������������������       �                      @        �       �                 ����?�q�q�?             @       �       �                    d@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   u@8�Z$���?             :@       �       �                   �Z@�8��8��?             8@        ������������������������       �                     �?        �       �                 ����?�nkK�?             7@        �       �                   �`@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        	             2@        ������������������������       �                      @        �       �                 ����?��۾%d�?#             M@       �       �                    b@�%^�?            �E@       �       �                   0a@�!���?             A@        ������������������������       �                     @        �       �                    �O@d��0u��?             >@        �       �                    �?     ��?             0@       �       �                   �`@�z�G��?             $@        ������������������������       �                     �?        �       �                    �N@�<ݚ�?             "@        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                   �^@և���X�?
             ,@       �       �                 ����?����X�?             @       �       �                   �j@      �?             @        ������������������������       �                     �?        �       �                   �p@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 `ff�?؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     "@        �       �                   �l@��S�ۿ?             .@        �       �                     P@      �?             @        ������������������������       �                      @        �       �                   �b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     &@        �                         �c@^�pӵL�?a            @d@       �                         �`@pJQg���?T            �`@       �       �                   �Q@(a��䛼?=            @Y@        �       �                    �N@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �                          �R@ ���v��?;            �X@       �       �                   pa@��8�$>�?9            @X@       ������������������������       �                    �J@        �       �                   �a@�C��2(�?             F@        �       �                   �]@�z�G��?             $@       ������������������������       �                     @        ������������������������       �                     @                               ����?г�wY;�?             A@                              ����?      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     :@                                p@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?              	                  `a@     ��?             @@        ������������������������       �                     @        
                        pl@ �Cc}�?             <@       ������������������������       �                     7@                                �b@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @                                  J@l��[B��?             =@                                �e@z�G�z�?             $@       ������������������������       �                     @                              ����?      �?             @        ������������������������       �                      @        ������������������������       �                      @                                 �?�����?             3@        ������������������������       �                     @                                 �?��
ц��?             *@                                �?�q�q�?             "@        ������������������������       �                     @                                 e@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KMKK��h^�B�   Np	�?���Gw{�?_���?B������?�{a���?5�rO#,�?�؉�؉�?�;�;�?)\���(�?�Q����?              �?l(�����?(������?UUUUUU�?UUUUUU�?              �?F]t�E�?]t�E]�?333333�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?�������?      �?                      �?      �?              �?              �?      �?F]t�E�?�.�袋�?UUUUUU�?UUUUUU�?              �?      �?                      �?333333�?ffffff�?UUUUUU�?UUUUUU�?              �?      �?        �$I�$I�?۶m۶m�?      �?      �?      �?                      �?              �?����?����?�$I�$I�?�m۶m��?333333�?333333�?333333�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?        _�_�?�A�A�?              �?333333�?�������?      �?                      �?�M1j���? Y����?              �?F]t�E�?]t�E]�?R���Q�?���Q��?ffffff�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?�������?�������?d!Y�B�?Nozӛ��?�������?�������?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?�؉�؉�?�;�;�?              �?�$I�$I�?۶m۶m�?۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?t�E]t�?F]t�E�?      �?      �?UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?                      �?�$I�$I�?۶m۶m�?              �?�������?�������?              �?      �?      �?      �?                      �?      �?        ۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?      �?                      �?      �?        
ףp=
�?=
ףp=�?�q�q�?��8��8�?      �?                      �?      �?      �?      �?      �?UUUUUU�?UUUUUU�?              �?      �?              �?        UUUUUU�?UUUUUU�?(�����?�5��P�?UUUUUU�?UUUUUU�?      �?                      �?              �?�������?�������?              �?      �?      �?      �?                      �?��h{��?�.�	��?��MbX�?9��v���?�)�B��?Y��~�?۬�ڬ��?�LɔL��?�F}g���?br1���?      �?      �?�$I�$I�?۶m۶m�?              �?      �?              �?        vb'vb'�?;�;��?333333�?�������?      �?        Cy�5��?^Cy�5�?�������?�������?�������?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?�������?�������?              �?UUUUUU�?UUUUUU�?              �?      �?              �?              �?        �|�ٓ�?a�2a�?E>�S��?�S�n�?)��?�[�w��?�������?�?ZZZZZZ�?�������?%I�$I��?�m۶m��?      �?              �?      �?              �?      �?        ffffff�?�������?      �?        �������?�������?      �?                      �?      �?              �?      �?�������?�������?      �?                      �?�m۶m��?�$I�$I�?      �?        �������?�������?      �?      �?��y��y�?�a�a�?      �?      �?      �?                      �?      �?        F]t�E�?/�袋.�?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?      �?        ��-��-�?�A�A�?      �?        UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?      �?      �?                      �?ؽ�u�{�?�E(B�?�B!��?���{��?�������?�������?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?        ;�;��?;�;��?UUUUUU�?UUUUUU�?      �?        d!Y�B�?�Mozӛ�?�������?�������?              �?      �?                      �?      �?        sO#,�4�?a����?�}A_��?�}A_�?�������?�������?      �?        DDDDDD�?wwwwww�?      �?      �?ffffff�?333333�?              �?9��8���?�q�q�?              �?      �?              �?        ۶m۶m�?�$I�$I�?�m۶m��?�$I�$I�?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        �$I�$I�?۶m۶m�?              �?      �?              �?        �?�������?      �?      �?              �?      �?      �?              �?      �?                      �?�<ݚ�?���Hx�?\�qA��?���7G��?�F�tj�?��~�X�?      �?      �?      �?                      �?1ogH�۩?�y;Cb�?����?�Q�/��?              �?F]t�E�?]t�E�?333333�?ffffff�?              �?      �?        �?�?      �?      �?              �?      �?                      �?      �?      �?              �?      �?              �?      �?      �?        ۶m۶m�?%I�$I��?              �?333333�?�������?      �?                      �?���=��?GX�i���?�������?�������?              �?      �?      �?      �?                      �?Q^Cy��?^Cy�5�?      �?        �;�;�?�؉�؉�?UUUUUU�?UUUUUU�?              �?333333�?�������?      �?                      �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJu�7hG        hNhG        hNhBKhDKhEh)h,K ��h.��R�(KK��h^�C              �?�t�bhQhchLC       ���R�hgKhhhkKh)h,K ��h.��R�(KK��hL�C       �t�bK��R�}�(hKhuM/hvh)h,K ��h.��R�(KM/��h}�B�K         �                 ����?p�Vv���?�           ��@                                ���ٿX~�pX��?�            �v@        ������������������������       �                     @               e                    @L@Zb��'��?�            `v@              \                    �?�q�q��?�             n@                                 �\@      �?}             i@                                  �l@8�A�0��?             6@              	                   �X@؇���X�?             ,@        ������������������������       �                     @        
                           �H@����X�?             @                                  �Z@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @                                   [@      �?              @       ������������������������       �                     @                                  @\@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?               +                    �D@��
}�?q            @f@                                  �c@�e�,��?"            �M@                                  �P@      �?              @       ������������������������       �                     @                                  �`@      �?             @        ������������������������       �                     �?        ������������������������       �                     @               *                   �b@������?            �I@              )                   `e@�����?            �H@              $                   Xq@X�Cc�?             <@                                 �o@�IєX�?             1@       ������������������������       �                     "@                #                   �a@      �?              @        !       "                   �p@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        %       (                   �a@"pc�
�?             &@        &       '                   p`@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     5@        ������������������������       �                      @        ,       [                   @g@����n�?O            �]@       -       R                   �b@p/3�d��?N            �]@       .       =                   �`@      �?(             N@       /       0                   �U@�ݜ�?            �C@        ������������������������       �                      @        1       :                 tff�?�L���?            �B@       2       3                   �b@�FVQ&�?            �@@       ������������������������       �                     :@        4       5                   �\@����X�?             @        ������������������������       �                     �?        6       9                   �g@r�q��?             @        7       8                   @_@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ;       <                    �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        >       A                    @G@�G��l��?             5@        ?       @                   0a@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        B       I                   �`@���Q��?             .@        C       D                    �G@���Q��?             @        ������������������������       �                     �?        E       H                    ^@      �?             @        F       G                    �I@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        J       O                    �J@�z�G��?             $@       K       N                    �I@���Q��?             @       L       M                   �m@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        P       Q                   �a@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        S       Z                    @H@XB���?&             M@       T       Y                    �?�FVQ&�?            �@@        U       X                   Pf@�<ݚ�?             "@        V       W                    d@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     8@        ������������������������       �                     9@        ������������������������       �                     �?        ]       b                   �q@      �?             D@       ^       _                   @Y@�X�<ݺ?             B@        ������������������������       �                     �?        `       a                 ����?��?^�k�?            �A@       ������������������������       �                     A@        ������������������������       �                     �?        c       d                   �`@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        f       �                   �a@vs�G��?M            �]@       g       �                    �R@C@Tu��?8            �U@       h       �                 833�?ҳ�wY;�?7            @U@       i       �                    �?l`N���?#            �J@       j                          �`@�L�lRT�?            �F@       k       p                   �W@��
ц��?             :@        l       o                   �l@r�q��?             @       m       n                   �[@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        q       x                    n@�G�z��?             4@       r       s                    @M@�q�q�?             (@        ������������������������       �                     @        t       u                    Y@      �?              @        ������������������������       �                      @        v       w                   �_@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        y       z                     N@      �?              @        ������������������������       �                      @        {       ~                   @_@      �?             @       |       }                   @`@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                   `d@�KM�]�?             3@       �       �                    a@r�q��?             (@        ������������������������       �                     @        �       �                    @N@�<ݚ�?             "@       �       �                    d@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �[@      �?              @        ������������������������       �                      @        ������������������������       �                     @        �       �                 ����?      �?             @@       �       �                   �a@��2(&�?             6@       �       �                    _@      �?	             0@        �       �                    ^@z�G�z�?             @        ������������������������       �                     @        �       �                   �o@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     &@        �       �                   @n@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                    �M@      �?             $@        ������������������������       �                     @        �       �                    �?r�q��?             @        ������������������������       �                     @        �       �                     O@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �d@�4�����?             ?@       �       �                    �N@�c�Α�?             =@        �       �                   �e@$�q-�?	             *@       ������������������������       �                     (@        ������������������������       �                     �?        �       �                   �a@     ��?             0@       �       �                   `c@      �?             (@        ������������������������       �                     @        �       �                    \@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �                          �?�zц��?�            w@       �                         �b@      �?�            @p@       �       �                 pff�?��r._�?�            �i@        �       �                 ����?r�qG�?A             X@       �       �                    �?�������?=            �U@       �       �                   �]@д>��C�?*             M@        �       �                   �s@���N8�?             5@       ������������������������       �                     4@        ������������������������       �                     �?        �       �                   �s@���"͏�?            �B@       �       �                   `a@�<ݚ�?             B@       �       �                   Hq@b�2�tk�?             2@       �       �                   �^@��
ц��?             *@        ������������������������       �                      @        �       �                   �`@���|���?
             &@        �       �                    �?r�q��?             @        ������������������������       �                      @        �       �                    �H@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?���Q��?             @       �       �                   �j@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                 033�?�X�<ݺ?             2@       ������������������������       �        	             .@        �       �                   �p@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   v@��>4և�?             <@       �       �                    �Q@$��m��?             :@       �       �                   �_@�q�q�?             8@       �       �                 033�?r�q��?             2@       �       �                    �L@8�Z$���?	             *@        �       �                   �Y@      �?             @        ������������������������       �                     �?        �       �                   @^@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     "@        �       �                   �^@z�G�z�?             @       �       �                    �N@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �a@�q�q�?             @        �       �                    �F@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        �       �                   @[@      �?             $@        ������������������������       �                     @        ������������������������       �                     @        �       �                    �J@��<nd�?D            @[@        �       �                   �Z@     ��?             @@        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    @J@\-��p�?             =@       �       �                    �D@`2U0*��?             9@        ������������������������       �                     �?        ������������������������       �                     8@        �       �                   �`@      �?             @       �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?`<)�+�?/            @S@        �       �                    `P@$�q-�?             :@       ������������������������       �                     3@        �       �                   �b@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        �                        `ff�?���J��?            �I@        �       �                    �?r�q��?             @        ������������������������       �                     @        �       �                   @l@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                    �F@                                Xr@�eP*L��?"            �K@                                �M@�q���?             H@                               �`@�q�q�?             B@                                �I@��Q��?             4@                                @B@��
ц��?	             *@        ������������������������       �                     @              	                   �B@�z�G��?             $@        ������������������������       �                     @        
                        �\@և���X�?             @                                pe@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?                                �e@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @                                `c@      �?	             0@                                 M@��S�ۿ?             .@       ������������������������       �                     &@                                �m@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?                                0n@r�q��?             (@                                �j@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @              $                  �k@��<nd�?N            @[@              !                033@�"w����?3             S@       ������������������������       �        0            @R@        "      #                   @O@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        %      (                   �J@r٣����?            �@@        &      '                  �p@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        )      .                   �N@؇���X�?             <@       *      -                  d@�<ݚ�?             2@       +      ,                   @N@      �?             0@       ������������������������       �                     ,@        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �        
             $@        �t�b��)     h�h)h,K ��h.��R�(KM/KK��h^�B�  w
��,@�?�z�����?�^�z���?�B�
*�?              �?x����X�?��¨N�?�������?UUUUUU�?      �?      �?/�袋.�?颋.���?�$I�$I�?۶m۶m�?              �?�$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?      �?      �?              �?      �?              �?      �?        ��d%+Y�?�MmjS��?�pR���?_[4��?      �?      �?              �?      �?      �?      �?                      �?xxxxxx�?�?^N��)x�?����X�?%I�$I��?�m۶m��?�?�?      �?              �?      �?      �?      �?              �?      �?              �?        F]t�E�?/�袋.�?      �?      �?              �?      �?                      �?      �?                      �?��(��(�?�\�\�?����c�?~ylE�p�?      �?      �?\��[���?�i�i�?              �?}���g�?L�Ϻ��?>����?|���?      �?        �m۶m��?�$I�$I�?              �?�������?UUUUUU�?      �?      �?              �?      �?              �?              �?      �?      �?                      �?1�0��?��y��y�?�������?UUUUUU�?              �?      �?        �������?333333�?333333�?�������?              �?      �?      �?      �?      �?      �?                      �?      �?        333333�?ffffff�?�������?333333�?      �?      �?      �?                      �?      �?        �������?�������?              �?      �?        GX�i���?�{a���?>����?|���?9��8���?�q�q�?333333�?�������?      �?                      �?      �?              �?              �?                      �?      �?      �?��8��8�?�q�q�?              �?_�_��?�A�A�?      �?                      �?      �?      �?              �?      �?        ���؊��?�N��?��C��:�?Ȥx�L��?�������?�������?�R���?
�[���?�I��I��?l�l��?�؉�؉�?�;�;�?UUUUUU�?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?�������?�������?UUUUUU�?UUUUUU�?      �?              �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?      �?              �?      �?      �?      �?      �?              �?      �?                      �?�k(���?(�����?�������?UUUUUU�?      �?        9��8���?�q�q�?      �?      �?      �?                      �?              �?      �?              �?      �?      �?                      �?      �?      �?��.���?t�E]t�?      �?      �?�������?�������?      �?              �?      �?              �?      �?              �?        UUUUUU�?UUUUUU�?      �?                      �?      �?      �?      �?        UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?��RJ)��?���Zk��?�{a���?5�rO#,�?;�;��?�؉�؉�?              �?      �?              �?      �?      �?      �?              �?333333�?�������?              �?      �?              �?              �?        o`E\��?@��(��?      �?      �?ە�]���?�ڕ�]��?UUUUUU�?UUUUUU�?��}A�?����/�?|a���?a���{�?�a�a�?��y��y�?              �?      �?        *�Y7�"�?v�)�Y7�?�q�q�?9��8���?9��8���?�8��8��?�;�;�?�؉�؉�?              �?]t�E]�?F]t�E�?�������?UUUUUU�?      �?              �?      �?              �?      �?        �������?333333�?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?�q�q�?��8��8�?              �?UUUUUU�?UUUUUU�?              �?      �?              �?        I�$I�$�?۶m۶m�?vb'vb'�?�N��N��?�������?�������?UUUUUU�?�������?;�;��?;�;��?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?�������?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?              �?              �?              �?              �?      �?              �?      �?        4R1�:#�?����[�?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?�{a���?a����?{�G�z�?���Q��?      �?                      �?      �?      �?      �?      �?              �?      �?              �?        ��O���?S{����?;�;��?�؉�؉�?              �?�$I�$I�?�m۶m��?              �?      �?        �?______�?UUUUUU�?�������?              �?      �?      �?              �?      �?                      �?t�E]t�?]t�E�?�������?�������?�������?�������?ffffff�?�������?�;�;�?�؉�؉�?              �?ffffff�?333333�?      �?        �$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?              �?      �?              �?      �?      �?                      �?              �?      �?      �?�������?�?      �?              �?      �?              �?      �?                      �?UUUUUU�?�������?�������?333333�?              �?      �?                      �?      �?        4R1�:#�?����[�?(�����?Cy�5��?              �?UUUUUU�?UUUUUU�?              �?      �?        |���?>���>�?�������?�������?      �?                      �?�$I�$I�?۶m۶m�?�q�q�?9��8���?      �?      �?              �?      �?              �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��!XhG        hNhG        hNhBKhDKhEh)h,K ��h.��R�(KK��h^�C              �?�t�bhQhchLC       ���R�hgKhhhkKh)h,K ��h.��R�(KK��hL�C       �t�bK��R�}�(hKhuM-hvh)h,K ��h.��R�(KM-��h}�B@K         �                   �`@U�ք�?�           ��@               '                   �e@�~6�]�?�            @u@               "                    `@�t`�4 �?N            �^@                                 �\@|�űN�?I            @]@                                  �Z@0�)AU��?$            �L@       ������������������������       �                     >@                                ����? 7���B�?             ;@                                   �?ףp=
�?             $@       	       
                    ]@r�q��?             @        ������������������������       �                     @                                   `@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     1@                                   �Q@�?�P�a�?%             N@                                  �?@4և���?"             L@       ������������������������       �                    �B@                                   п���y4F�?             3@        ������������������������       �                     �?                                  �]@r�q��?
             2@        ������������������������       �                     @                                    P@���!pc�?             &@                                  @O@և���X�?             @                                  `@z�G�z�?             @        ������������������������       �                     @                                  �`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @                !                 ����?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        #       $                 ����?���Q��?             @        ������������������������       �                      @        %       &                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        (                          p`@"wO�a��?�            @k@       )       `                   �`@�WV�?�             j@        *       [                    �?��9܂�?=            @V@       +       N                    �?a��t��?7            �S@       ,       7                   �j@V{q֛w�?+             O@        -       2                 @33�?��Q��?             4@        .       1                    @H@����X�?             @        /       0                   �]@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        3       6                   �h@8�Z$���?             *@       4       5                    �G@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        8       ?                   0o@�q�q�?             E@        9       >                    �?��s����?             5@        :       ;                   �k@z�G�z�?             @        ������������������������       �                      @        <       =                   �l@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �        	             0@        @       M                 ����?�G��l��?             5@       A       F                 ����?      �?             0@        B       E                   hs@X�<ݚ�?             "@       C       D                     N@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        G       H                 433�?����X�?             @        ������������������������       �                     �?        I       L                   Hr@�q�q�?             @        J       K                   Hq@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        O       Z                    `@      �?             0@       P       S                   @Z@����X�?
             ,@        Q       R                    �K@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        T       U                   �k@�����H�?             "@        ������������������������       �                     @        V       Y                    @M@r�q��?             @        W       X                   �_@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        \       ]                   �g@"pc�
�?             &@        ������������������������       �                     �?        ^       _                   �T@ףp=
�?             $@        ������������������������       �                     �?        ������������������������       �                     "@        a       x                    �?�p�I�?H            �]@       b       o                 `ff�?p�}�ޤ�?/            @R@        c       d                    �?���y4F�?             3@        ������������������������       �                      @        e       n                   �a@�t����?             1@       f       m                    �P@z�G�z�?             $@       g       l                    �L@�����H�?             "@        h       k                    _@      �?             @       i       j                 hff�?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        p       u                   @s@�>����?!             K@       q       r                 `ff@ qP��B�?            �E@       ������������������������       �                     C@        s       t                 ���@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        v       w                    �Q@���!pc�?             &@       ������������������������       �                      @        ������������������������       �                     @        y       ~                 ����?���.�6�?             G@        z       {                   �h@�θ�?             *@        ������������������������       �                      @        |       }                    �I@�C��2(�?             &@        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                    �@@        ������������������������       �                     $@        �       �                    @L@�����?           �x@       �       �                    �?6通(��?�            �p@       �       �                   @W@���0��?�            �m@        ������������������������       �                     @        �       �                   @E@���2���?�            `m@        ������������������������       �                      @        �       �                 033@8ӈ(�3�?�             m@       �       �                 ����?&^�r���?�            @l@       �       �                    @C@x�ۈp�?u            `e@        �       �                   �f@���N8�?             5@       �       �                   �c@X�Cc�?             ,@        ������������������������       �                      @        �       �                    �B@      �?             (@       ������������������������       �                      @        �       �                   0g@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                   �g@ףp=
�?e            �b@       �       �                   a@��7*��?d            �b@        �       �                   �`@����X�?             @        ������������������������       �                     @        �       �                   0a@      �?             @        ������������������������       �                     �?        �       �                    @J@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                   �o@@�j;��?]            �a@       �       �                    @D@ p�/��?9            @V@        �       �                   `k@r�q��?             @        ������������������������       �                     @        �       �                   �l@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   k@P��BNֱ?5            �T@       �       �                   �j@��(\���?             D@       �       �                    �E@�7��?            �C@        ������������������������       �                     &@        �       �                    �?@4և���?             <@        �       �                   �e@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �b@ ��WV�?             :@       ������������������������       �        
             .@        �       �                   g@�C��2(�?             &@        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                     �?        ������������������������       �                    �E@        �       �                    �?f1r��g�?$            �J@        �       �                    ^@$�q-�?             *@        �       �                   �[@      �?             @        ������������������������       �                      @        �       �                    @E@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        �       �                   �e@z�G�z�?             D@       �       �                   0d@4?,R��?             B@       �       �                     E@      �?             4@        ������������������������       �                     @        �       �                    �J@X�Cc�?             ,@       �       �                   pa@      �?              @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     0@        �       �                   �q@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    @C@���!pc�?&            �K@        ������������������������       �                      @        �       �                    �G@�c�����?$            �J@        ������������������������       �                     0@        �       �                    �I@^H���+�?            �B@       �       �                 ����?      �?             4@       �       �                   �`@X�Cc�?             ,@       �       �                   �\@����X�?             @        ������������������������       �                     �?        �       �                 ����?r�q��?             @        �       �                    �H@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?r�q��?             @       �       �                   �`@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?@�0�!��?
             1@       ������������������������       �                     (@        �       �                   @b@���Q��?             @       �       �                    �J@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   g@����X�?             @       �       �                    \@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                    _@�4�����?             ?@        �       �                    �G@�q�q�?             (@        ������������������������       �                     @        ������������������������       �                     @        �       �                   �`@�S����?             3@       ������������������������       �                     &@        �       �                    �?      �?              @       �       �                    �?����X�?             @        �       �                    d@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �       �                   Pa@z�m�(�?N            @_@        �       �                   m@r�q��?             (@        �       �                    @N@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �                         pl@��\20�?F            @\@        �                         �O@v ��?            �E@        �       �                   �a@     ��?
             0@        ������������������������       �                      @        �                           `@@4և���?	             ,@       ������������������������       �                     $@                                �c@      �?             @       ������������������������       �                     @        ������������������������       �                     �?              	                  `b@��}*_��?             ;@                              `ff�?�n_Y�K�?
             *@                                �?����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        
                        �b@؇���X�?
             ,@                               Pe@      �?              @                               �i@؇���X�?             @                                 �M@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @              "                `ff�?���L��?(            �Q@              !                ����?��
ц��?             :@                              ����?
;&����?             7@                               Xr@b�2�tk�?
             2@                                 @O@"pc�
�?             &@                                �c@�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @                                 �?����X�?             @        ������������������������       �                     @                                @`@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        #      (                   �?t��ճC�?             F@       $      %                  �b@�X�<ݺ?             B@       ������������������������       �                     6@        &      '                   @P@؇���X�?             ,@       ������������������������       �                     (@        ������������������������       �                      @        )      *                   d@      �?              @        ������������������������       �                     @        +      ,                  �q@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �t�bh�h)h,K ��h.��R�(KM-KK��h^�B�  ᓔ��?�5�;��?�?999999�?�����?~�K�`�?���?�������?p�}��?��Gp�?              �?h/�����?	�%����?�������?�������?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?�����ݽ?DDDDDD�?�$I�$I�?n۶m۶�?              �?(������?6��P^C�?      �?        UUUUUU�?�������?              �?t�E]t�?F]t�E�?۶m۶m�?�$I�$I�?�������?�������?              �?      �?      �?      �?                      �?      �?                      �?      �?      �?              �?      �?        333333�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?        �߅���?�p=��?O��N���?ى�؉��?�.p��? ��G?��?��[��[�?!� ��?�{����?B!��?�������?ffffff�?�$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?              �?      �?                      �?;�;��?;�;��?�m۶m��?�$I�$I�?              �?      �?              �?        UUUUUU�?UUUUUU�?�a�a�?z��y���?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?��y��y�?1�0��?      �?      �?r�q��?�q�q�?�m۶m��?�$I�$I�?      �?                      �?              �?�m۶m��?�$I�$I�?      �?        UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?      �?      �?�m۶m��?�$I�$I�?�������?333333�?              �?      �?        �q�q�?�q�q�?      �?        �������?UUUUUU�?      �?      �?      �?                      �?      �?                      �?F]t�E�?/�袋.�?      �?        �������?�������?      �?                      �?���?:�:��?�
*T��?�z��ի�?6��P^C�?(������?              �?<<<<<<�?�?�������?�������?�q�q�?�q�q�?      �?      �?      �?      �?              �?      �?              �?              �?                      �?      �?        h/�����?�Kh/��?�}A_З?��}A�?              �?�������?�������?      �?                      �?t�E]t�?F]t�E�?              �?      �?        Y�B��?���7���?�؉�؉�?ى�؉��?      �?        F]t�E�?]t�E�?      �?                      �?              �?              �?R��3�M�?\e
�d�?%�N!&�?l�z�g�?����?X�3X�3�?              �?2���G�?�7'�h��?              �?/�祁�?C˯`h��?=���S�?+=����?�w�A�?�A|�?�a�a�?��y��y�?%I�$I��?�m۶m��?              �?      �?      �?      �?              �?      �?      �?                      �?      �?        �������?�������?]"<)H��?����?�m۶m��?�$I�$I�?      �?              �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?w�'�K�?H���@��?�G?�я�?p�\��?�������?UUUUUU�?      �?              �?      �?              �?      �?        ��FS���?���ˊ��?�������?333333�?��[��[�?�A�A�?      �?        n۶m۶�?�$I�$I�?      �?      �?      �?                      �?O��N���?;�;��?      �?        ]t�E�?F]t�E�?              �?      �?                      �?      �?        �!5�x+�?�x+�R�?�؉�؉�?;�;��?      �?      �?      �?              �?      �?      �?                      �?      �?        ffffff�?ffffff�?�8��8��?r�q��?      �?      �?      �?        %I�$I��?�m۶m��?      �?      �?      �?                      �?      �?              �?              �?      �?              �?      �?                      �?F]t�E�?t�E]t�?              �?�V�9�&�?:�&oe�?      �?        L�Ϻ��?�g�`�|�?      �?      �?�m۶m��?%I�$I��?�m۶m��?�$I�$I�?              �?�������?UUUUUU�?      �?      �?              �?      �?              �?                      �?�������?UUUUUU�?�������?�������?      �?                      �?      �?        ZZZZZZ�?�������?      �?        �������?333333�?UUUUUU�?UUUUUU�?      �?                      �?              �?�$I�$I�?�m۶m��?UUUUUU�?�������?      �?                      �?      �?        ��RJ)��?���Zk��?�������?�������?              �?      �?        ^Cy�5�?(������?              �?      �?      �?�$I�$I�?�m۶m��?      �?      �?              �?      �?                      �?      �?        ���Mb�?+�����?�������?UUUUUU�?333333�?�������?              �?      �?              �?        �JO-���?�ZX驅�?qG�w��?G�w��?      �?      �?      �?        �$I�$I�?n۶m۶�?              �?      �?      �?              �?      �?        _B{	�%�?B{	�%��?ى�؉��?;�;��?�m۶m��?�$I�$I�?      �?                      �?              �?۶m۶m�?�$I�$I�?      �?      �?۶m۶m�?�$I�$I�?      �?      �?      �?                      �?      �?                      �?      �?        _�_��?��:��:�?�;�;�?�؉�؉�?�Mozӛ�?Y�B��?�8��8��?9��8���?/�袋.�?F]t�E�?UUUUUU�?UUUUUU�?      �?                      �?      �?        �$I�$I�?�m۶m��?              �?      �?      �?      �?                      �?              �?      �?        t�E]t�?�E]t��?�q�q�?��8��8�?              �?�$I�$I�?۶m۶m�?              �?      �?              �?      �?              �?      �?      �?              �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJC�NhG        hNhG        hNhBKhDKhEh)h,K ��h.��R�(KK��h^�C              �?�t�bhQhchLC       ���R�hgKhhhkKh)h,K ��h.��R�(KK��hL�C       �t�bK��R�}�(hKhuMOhvh)h,K ��h.��R�(KMO��h}�B�S         �                 ����?4�5����?�           ��@                                 @E@�Ff��K�?�            x@                                  �[@��x_F-�?#            �I@        ������������������������       �                     3@                                  �]@     ��?             @@                                   @N@X�<ݚ�?             "@                                  @\@z�G�z�?             @        ������������������������       �                      @        	       
                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                   �?      �?             @                                  �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @                                   @O@��<b���?             7@                                  a@�KM�]�?             3@        ������������������������       �                     $@                                   \@�<ݚ�?             "@                                  `b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                   �?؇���X�?             @                                hff�?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @                                ����?      �?             @        ������������������������       �                     �?        ������������������������       �                     @                �                 ����?:�{��x�?�            �t@       !       R                   `_@&���(�?�            �s@        "       K                   �p@������?-            @Q@       #       J                 hff�?l��[B��?&             M@       $       %                    �F@�eP*L��?$            �K@        ������������������������       �                     @        &       I                     P@���Q��?"             I@       '       (                   �V@\X��t�?             G@        ������������������������       �                     @        )       H                   �^@�ՙ/�?             E@       *       C                    @M@X�<ݚ�?             B@       +       ,                   �d@��>4և�?             <@        ������������������������       �                      @        -       B                    �?$��m��?             :@       .       /                    @H@և���X�?             5@        ������������������������       �                      @        0       A                   o@p�ݯ��?             3@       1       <                    �?�q�q�?             2@       2       ;                    ^@������?             .@       3       8                   �l@d}h���?             ,@       4       7                    Z@      �?              @        5       6                    @J@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        9       :                    �J@�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        =       >                     K@�q�q�?             @        ������������������������       �                     �?        ?       @                   �\@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        D       E                   @k@      �?              @        ������������������������       �                     @        F       G                    �O@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        L       M                   �q@"pc�
�?             &@       ������������������������       �                      @        N       O                   �r@�q�q�?             @        ������������������������       �                     �?        P       Q                   @[@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        S       h                    �?^�pӵL�?�            `n@        T       U                   �[@`�Q��?$             I@        ������������������������       �                     @        V       g                   �d@��+7��?"             G@       W       Z                   �_@RB)��.�?             �E@        X       Y                   Xq@X�Cc�?	             ,@       ������������������������       �                     "@        ������������������������       �                     @        [       b                   �b@\-��p�?             =@        \       ]                    �H@�q�q�?             "@        ������������������������       �                     �?        ^       _                   �?      �?              @       ������������������������       �                     @        `       a                    �K@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        c       d                    �M@P���Q�?             4@       ������������������������       �                     ,@        e       f                   8r@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        i       �                   �t@��y�S��?{             h@       j       s                   Pg@��r
'��?w            @g@        k       p                   ``@��a�n`�?             ?@       l       o                    �?�q�q�?
             2@       m       n                   �f@؇���X�?	             ,@       ������������������������       �                     (@        ������������������������       �                      @        ������������������������       �                     @        q       r                   f@$�q-�?	             *@       ������������������������       �                     (@        ������������������������       �                     �?        t       �                    �P@(�����?d            `c@       u       �                    c@�:�]��?b             c@        v       �                   �[@��ɉ�?*            @P@        w       |                   @[@      �?	             0@       x       {                 ����?�����H�?             "@       y       z                    m@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        }       ~                   `a@����X�?             @        ������������������������       �                     �?               �                   �a@r�q��?             @        ������������������������       �                     @        �       �                    @G@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �d@��<D�m�?!            �H@       �       �                    �H@ �q�q�?              H@        ������������������������       �                     9@        �       �                 ����?���}<S�?             7@       �       �                   �b@�r����?             .@       �       �                   �k@$�q-�?	             *@        �       �                   �j@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   0a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                    b@�zvܰ?8             V@       �       �                   �e@ �й���?0            @R@       ������������������������       �        $             K@        �       �                   @p@�}�+r��?             3@       ������������������������       �                     2@        ������������������������       �                     �?        �       �                    @L@�r����?             .@       �       �                   �f@�8��8��?             (@       ������������������������       �                     &@        ������������������������       �                     �?        �       �                   �d@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   `c@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?؇���X�?             @       �       �                    `@      �?             @        ������������������������       �                     �?        �       �                    �J@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?�eP*L��?
             6@       �       �                    �?      �?	             0@        �       �                   �c@      �?              @       �       �                   �q@r�q��?             @       �       �                   �`@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        �       �                    @I@      �?              @       �       �                    �H@���Q��?             @       ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �                         �`@�?ʵ���?�            �u@       �       �                 pff�?���U��?z            @g@       �       �                   0b@�X���?H             \@        �       �                    @K@�g�y��?             ?@        �       �                    @J@@4և���?
             ,@       ������������������������       �                     (@        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        
             1@        �       �                   Xy@LMc����?4            @T@       �       �                    �D@J�����?2            @S@        �       �                   e@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        �       �                   �t@�l�]�N�?,             Q@       �       �                   @Z@���Q��?)            @P@        ������������������������       �                     @        �       �                   `W@��Q��?&             N@        ������������������������       �                     @        �       �                   �e@Dc}h��?$             L@       �       �                     M@�q�q�?"            �I@       �       �                 ����?��Q���?             D@       �       �                    `@8�A�0��?             6@       �       �                    _@      �?	             (@       �       �                   0m@���Q��?             $@        �       �                    �I@���Q��?             @       �       �                     G@      �?             @       �       �                   ``@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �p@z�G�z�?             @        ������������������������       �                     @        �       �                   `]@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �`@�z�G��?             $@       �       �                    �?�q�q�?             "@        �       �                   �]@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �j@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    \@�����H�?
             2@        ������������������������       �                     �?        �       �                    �J@�IєX�?	             1@       ������������������������       �                     "@        �       �                    �?      �?              @        ������������������������       �                     @        �       �                   @a@      �?             @        ������������������������       �                     �?        �       �                   �o@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �k@�eP*L��?
             &@        ������������������������       �                      @        �       �                   �p@�q�q�?             "@        ������������������������       �                     @        �       �                   xr@      �?             @        ������������������������       �                      @        �       �                   �`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @                                  �F@�x
�2�?2            �R@                                @_@X�<ݚ�?             "@                                �?r�q��?             @                                �`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @                                 _@ ����?+            @P@        	                        `l@z�G�z�?             >@        
                         @N@X�Cc�?	             ,@                               `U@      �?              @                               @^@      �?             @                             ��� @      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @                                @]@      �?             0@                                pp@z�G�z�?             @                              ���@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     &@                                  O@��?^�k�?            �A@       ������������������������       �                     <@                                 �?؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?              @                  �b@D���\�?p            `d@              )                  0`@@4և���?\            �a@       !      &                   �Q@��'cy�??            @Y@       "      %                  `l@�L��ȕ?;            @W@       #      $                  0l@��<b�ƥ?             G@       ������������������������       �                    �F@        ������������������������       �                     �?        ������������������������       �                    �G@        '      (                  �c@      �?              @        ������������������������       �                     @        ������������������������       �                     @        *      3                   @K@8�Z$���?            �C@        +      ,                   @J@����X�?
             ,@        ������������������������       �                     @        -      .                   �?      �?              @        ������������������������       �                      @        /      2                   �?�q�q�?             @       0      1                   �J@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        4      7                  �N@HP�s��?             9@        5      6                    N@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        8      ?                  `a@���7�?             6@        9      >                   �?      �?              @       :      ;                  �b@      �?             @        ������������������������       �                      @        <      =                   @Q@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     ,@        A      N                   e@�û��|�?             7@       B      M                `ff@և���X�?             5@       C      D                  `c@��.k���?             1@        ������������������������       �                     @        E      F                   @F@և���X�?             ,@        ������������������������       �                      @        G      L                  �d@�q�q�?             (@       H      K                  �c@      �?              @       I      J                  �r@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �t�bh�h)h,K ��h.��R�(KMOKK��h^�B�   Np	�?���Gw{�?��2�q�?��?�?�������?              �?      �?      �?r�q��?�q�q�?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?      �?      �?      �?              �?      �?                      �?��Moz��?��,d!�?(�����?�k(���?              �?�q�q�?9��8���?      �?      �?      �?                      �?�$I�$I�?۶m۶m�?      �?      �?      �?                      �?              �?      �?      �?              �?      �?        �R&����?qZ�}�z�?�i�i�?��[��[�??���(�?ہ�v`��?GX�i���?���=��?]t�E�?t�E]t�?      �?        �������?333333�?��Moz��?!Y�B�?      �?        �a�a�?�<��<��?�q�q�?r�q��?I�$I�$�?۶m۶m�?      �?        vb'vb'�?�N��N��?۶m۶m�?�$I�$I�?      �?        Cy�5��?^Cy�5�?UUUUUU�?UUUUUU�?�?wwwwww�?۶m۶m�?I�$I�$�?      �?      �?      �?      �?              �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?              �?        UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?      �?                      �?      �?      �?      �?              �?      �?              �?      �?                      �?              �?      �?        /�袋.�?F]t�E�?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?        ���Hx�?�<ݚ�?��(\���?{�G�z�?              �?zӛ����?Y�B��?S֔5eM�?���)k��?%I�$I��?�m۶m��?      �?                      �?a����?�{a���?UUUUUU�?UUUUUU�?              �?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?ffffff�?�������?      �?        �������?UUUUUU�?      �?                      �?              �?�l.j��?�LF�W>�?�<��#��?�n�ᆻ?�c�1��?�s�9��?UUUUUU�?UUUUUU�?۶m۶m�?�$I�$I�?      �?                      �?              �?�؉�؉�?;�;��?      �?                      �?Q���P�?y�W�x�?}}}}}}�?�?�����?�����?      �?      �?�q�q�?�q�q�?�������?�������?      �?                      �?      �?        �$I�$I�?�m۶m��?      �?        UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?              �?      �?        ��S�r
�?և���X�?�������?UUUUUU�?      �?        ӛ���7�?d!Y�B�?�������?�?�؉�؉�?;�;��?�������?�������?      �?                      �?      �?              �?      �?      �?                      �?      �?                      �?颋.���?t�E]t�?����Ǐ�?����?      �?        �5��P�?(�����?      �?                      �?�������?�?UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?              �?      �?              �?      �?        �$I�$I�?۶m۶m�?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?]t�E�?t�E]t�?      �?      �?      �?      �?�������?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?      �?      �?�������?333333�?      �?                      �?      �?                      �?`�tՁ�?��ע��?EM4�D�?^v�e�]�?n۶m۶�?I�$I�$�?�B!��?��{���?�$I�$I�?n۶m۶�?              �?      �?      �?              �?      �?                      �?��ӭ�a�?k~X�<�?V~B����?S{����?�q�q�?�q�q�?              �?      �?        ZZZZZZ�?KKKKKK�?333333�?�������?              �?�������?ffffff�?              �?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?333333�?�������?颋.���?/�袋.�?      �?      �?333333�?�������?�������?333333�?      �?      �?      �?      �?              �?      �?                      �?      �?        �������?�������?      �?              �?      �?      �?                      �?              �?ffffff�?333333�?UUUUUU�?UUUUUU�?      �?      �?              �?      �?        333333�?�������?      �?                      �?      �?        �q�q�?�q�q�?              �?�?�?      �?              �?      �?      �?              �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?        ]t�E�?t�E]t�?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?      �?              �?      �?      �?                      �?      �?                      �?      �?        o0E>��?�n0E>�?�q�q�?r�q��?UUUUUU�?�������?      �?      �?              �?      �?                      �?      �?        �����?�ȍ�ȍ�?�������?�������?�m۶m��?%I�$I��?      �?      �?      �?      �?      �?      �?      �?                      �?              �?      �?                      �?      �?      �?�������?�������?      �?      �?              �?      �?                      �?              �?�A�A�?_�_��?              �?�$I�$I�?۶m۶m�?              �?      �?        ��g*׽?n�
�E�?�$I�$I�?n۶m۶�?��be�F�?`ҩy���?X`��?��~���?d!Y�B�?��7��M�?              �?      �?                      �?      �?      �?              �?      �?        ;�;��?;�;��?�$I�$I�?�m۶m��?              �?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?                      �?              �?{�G�z�?q=
ףp�?UUUUUU�?UUUUUU�?      �?                      �?F]t�E�?�.�袋�?      �?      �?      �?      �?              �?      �?      �?      �?                      �?              �?              �?��,d!�?8��Moz�?۶m۶m�?�$I�$I�?�������?�?      �?        ۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?      �?      �?�������?�������?              �?      �?              �?                      �?              �?              �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�R�[hG        hNhG        hNhBKhDKhEh)h,K ��h.��R�(KK��h^�C              �?�t�bhQhchLC       ���R�hgKhhhkKh)h,K ��h.��R�(KK��hL�C       �t�bK��R�}�(hKhuM1hvh)h,K ��h.��R�(KM1��h}�B@L         �                   �a@6������?�           ��@              �                    �?�" ED��?f           ��@                                 �_@��It��?�            �s@                                   @D@�����?            �H@        ������������������������       �                      @                                  P`@���?            �D@                                  \@z�G�z�?             >@                                   `@�q�q�?             "@       	                           �?r�q��?             @       
                          @\@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @                                   d@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?                                   �?؇���X�?             5@                                 �`@$�q-�?	             *@       ������������������������       �                     (@        ������������������������       �                     �?                                  �\@      �?              @       ������������������������       �                     @        ������������������������       �                      @                                ����?���|���?             &@        ������������������������       �                     @                                   �?z�G�z�?             @                                  �N@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?               ~                    �Q@�+���-�?�            �p@               Y                    @L@@�4���?�            Pp@       !       ,                   a@|�%�9��?�             i@        "       +                   r@">�֕�?            �A@       #       $                    �F@z�G�z�?             >@        ������������������������       �                     "@        %       &                   �]@����X�?             5@        ������������������������       �                     @        '       (                    �J@      �?
             0@       ������������������������       �                      @        )       *                   a@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        -       @                   0n@��Lɿ��?k            �d@       .       5                    �D@�nkK�?=             W@        /       4                   �d@�����H�?             ;@        0       3                   �\@�z�G��?             $@        1       2                   @c@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �        
             1@        6       ?                   Pi@ ����?+            @P@        7       8                   �b@ �q�q�?             8@        ������������������������       �                     $@        9       >                   �c@@4և���?	             ,@        :       ;                     F@r�q��?             @        ������������������������       �                     @        <       =                   @_@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                    �D@        A       V                 ����?��G���?.            �R@       B       I                   `]@��a�2��?,             R@        C       H                    �H@      �?
             4@       D       G                     G@�θ�?             *@       E       F                    q@      �?              @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        J       K                   `_@0G���ջ?"             J@        ������������������������       �                     .@        L       Q                    �?�L���?            �B@       M       P                    �B@�g�y��?             ?@        N       O                     @@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     ;@        R       S                    @I@�q�q�?             @        ������������������������       �                     �?        T       U                   0`@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        W       X                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        Z       s                    @N@      �?)             N@       [       r                   Ps@X�Cc�?             <@       \       m                   ``@���Q��?             9@       ]       b                    �?���Q��?             .@        ^       a                 ����?r�q��?             @        _       `                    �L@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        c       l                 ����?X�<ݚ�?             "@       d       e                   @Z@և���X�?             @        ������������������������       �                     �?        f       g                   �f@�q�q�?             @        ������������������������       �                     �?        h       i                   �_@z�G�z�?             @        ������������������������       �                      @        j       k                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        n       q                   @f@ףp=
�?             $@        o       p                   �b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        t       }                    �?     ��?             @@       u       x                    �?���B���?             :@        v       w                   `V@      �?             @        ������������������������       �                     @        ������������������������       �                     @        y       |                    �?ףp=
�?             4@       z       {                   @t@"pc�
�?             &@       ������������������������       �                     "@        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                     @               �                    �?r�q��?             @       �       �                 ����?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?4ӏEI�?�            `o@       �       �                   Pg@����X�?}            `i@        �       �                   �_@���c���?             J@        �       �                    @p�ݯ��?             3@       �       �                 ����?      �?
             ,@        �       �                   pf@      �?              @       �       �                    I@����X�?             @        �       �                   �O@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �       �                   @^@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                    �@@        �       �                    �L@�� �\��?^            �b@       �       �                    �A@��MΖ��?:            @W@        ������������������������       �                     @        �       �                 033�?������?7            �U@       �       �                   �[@j���� �?             �I@        �       �                 ����?�z�G��?             $@       �       �                 ����?      �?              @       �       �                    b@؇���X�?             @        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �J@#z�i��?            �D@       �       �                    �G@�eP*L��?             6@        �       �                    �?"pc�
�?             &@       �       �                   �b@ףp=
�?             $@        �       �                   �m@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?���!pc�?	             &@        ������������������������       �                     �?        �       �                    a@z�G�z�?             $@       �       �                 ����?����X�?             @        ������������������������       �                     �?        �       �                 ����?r�q��?             @        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                   8t@���y4F�?
             3@       �       �                   �_@�t����?             1@       �       �                   �g@z�G�z�?             $@        ������������������������       �                     �?        �       �                 ����?�����H�?             "@       ������������������������       �                     @        �       �                   b@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        �       �                 ���@*O���?             B@       �       �                   pp@h+�v:�?             A@       �       �                   b@
;&����?             7@       �       �                    @������?	             .@       �       �                   �`@ףp=
�?             $@       ������������������������       �                      @        �       �                   �j@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    n@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        �       �                     I@�C��2(�?             &@        �       �                    @�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        �       �                     R@\-��p�?$             M@       �       �                   �h@���5��?#            �L@        ������������������������       �                     �?        �       �                   �a@ �Cc}�?"             L@       �       �                    ^@      �?             @@        �       �                    �N@@4և���?             ,@        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     (@        ������������������������       �                     2@        �       �                    @�q�q�?             8@       �       �                    �?�t����?
             1@        �       �                   �\@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �c@      �?              @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?8��8���?             H@        �       �                   �a@      �?             @       ������������������������       �                      @        ������������������������       �                      @        �       �                   �x@t��ճC�?             F@       �       �                   �c@�Ń��̧?             E@       ������������������������       �                     B@        �       �                    �I@r�q��?             @        ������������������������       �                     @        �       �                 `ff@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       $                pff�?L�e[���?g            �d@       �       �                   �b@bOvj6��?E            �[@        �       �                    �?��2(&�?             6@        �       �                   �a@      �?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �        	             0@        �       �                   @\@~�4_�g�?9             V@        ������������������������       �                     0@                                 @]@)O���?-             R@                                `c@�����H�?             "@                                 @K@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @                                ph@�G��l��?(            �O@                                 �?��s����?             5@       ������������������������       �                     $@        	                      ����?���|���?             &@       
                        �c@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @                                `k@�ՙ/�?             E@        ������������������������       �                      @                                 s@��.k���?             A@                                �?�q�q�?             8@                               �_@������?             1@        ������������������������       �                     @                                 �B@���|���?             &@        ������������������������       �                     �?                                �n@�z�G��?             $@                                 F@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @                                pd@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?              #                   �?z�G�z�?             $@             "                   �?�����H�?             "@               !                ����?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        %      (                   �?�}�+r��?"            �L@        &      '                   @P@      �?	             0@       ������������������������       �                     ,@        ������������������������       �                      @        )      *                `ff@��Y��]�?            �D@       ������������������������       �                     <@        +      0                   �?$�q-�?	             *@       ,      /                  �l@�����H�?             "@        -      .                  @c@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �t�b��     h�h)h,K ��h.��R�(KM1KK��h^�B  ��X�5�?��S�$e�?�\l�?t���G'�?-n����?�#{���?����X�?^N��)x�?              �?8��18�?28��1�?�������?�������?UUUUUU�?UUUUUU�?UUUUUU�?�������?      �?      �?      �?                      �?              �?UUUUUU�?UUUUUU�?      �?                      �?�$I�$I�?۶m۶m�?;�;��?�؉�؉�?              �?      �?              �?      �?              �?      �?        F]t�E�?]t�E]�?              �?�������?�������?      �?      �?              �?      �?              �?        �e�h� �?xi�]�}�?=ZT"���?��v��?�N��b�?$�6��w�?_�_��?�A�A�?�������?�������?      �?        �m۶m��?�$I�$I�?              �?      �?      �?      �?              �?      �?      �?                      �?              �?�������?rY1P»?�Mozӛ�?d!Y�B�?�q�q�?�q�q�?ffffff�?333333�?      �?      �?      �?                      �?      �?              �?         �����? �����?�������?UUUUUU�?      �?        n۶m۶�?�$I�$I�?�������?UUUUUU�?      �?              �?      �?              �?      �?              �?              �?        #�u�)��?v�)�Y7�?��8��8�?�q�q�?      �?      �?�؉�؉�?ى�؉��?      �?      �?      �?                      �?              �?      �?        vb'vb'�?�؉�؉�?      �?        }���g�?L�Ϻ��?��{���?�B!��?      �?      �?      �?                      �?      �?        UUUUUU�?UUUUUU�?              �?�������?�������?              �?      �?              �?      �?              �?      �?              �?      �?%I�$I��?�m۶m��?333333�?�������?�������?333333�?UUUUUU�?�������?      �?      �?      �?                      �?              �?r�q��?�q�q�?۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?      �?        �������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        �������?�������?      �?      �?      �?                      �?      �?              �?              �?      �?��؉���?ى�؉��?      �?      �?      �?                      �?�������?�������?/�袋.�?F]t�E�?      �?                      �?      �?              �?        UUUUUU�?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?4���Q�?f4���?�$I�$I�?�m۶m��?�;�;�?;�;��?Cy�5��?^Cy�5�?      �?      �?      �?      �?�$I�$I�?�m۶m��?      �?      �?              �?      �?                      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?              �?�vV;���?��Tb*1�?�]v�e��?4�DM4�?              �?m��֡�?J��/�?�������?ZZZZZZ�?333333�?ffffff�?      �?      �?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?      �?        �+Q��?ە�]���?t�E]t�?]t�E�?/�袋.�?F]t�E�?�������?�������?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?t�E]t�?F]t�E�?      �?        �������?�������?�$I�$I�?�m۶m��?      �?        UUUUUU�?�������?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?6��P^C�?(������?<<<<<<�?�?�������?�������?              �?�q�q�?�q�q�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?                      �?�q�q�?�q�q�?xxxxxx�?�������?Y�B��?�Mozӛ�?�?wwwwww�?�������?�������?              �?      �?      �?              �?      �?        333333�?�������?              �?      �?              �?        F]t�E�?]t�E�?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?�{a���?a����?��Gp�?�}��?      �?        ۶m۶m�?%I�$I��?      �?      �?�$I�$I�?n۶m۶�?      �?      �?      �?                      �?              �?              �?�������?UUUUUU�?�������?�������?�q�q�?�q�q�?      �?                      �?      �?      �?      �?                      �?              �?      �?        �������?�������?      �?      �?              �?      �?        t�E]t�?�E]t��?�a�a�?��<��<�?              �?UUUUUU�?�������?              �?      �?      �?      �?                      �?      �?        3	v���?g�D����?�7�}���?�)A��?t�E]t�?��.���?      �?      �?      �?                      �?              �?��.���?/�袋.�?              �?9��8���?��8��8�?�q�q�?�q�q�?      �?      �?      �?                      �?      �?        ��y��y�?1�0��?�a�a�?z��y���?              �?F]t�E�?]t�E]�?      �?      �?      �?                      �?      �?        �<��<��?�a�a�?      �?        �������?�?�������?�������?�?xxxxxx�?              �?F]t�E�?]t�E]�?      �?        333333�?ffffff�?333333�?�������?              �?      �?                      �?۶m۶m�?�$I�$I�?      �?                      �?�������?�������?�q�q�?�q�q�?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?(�����?�5��P�?      �?      �?              �?      �?        ������?8��18�?              �?;�;��?�؉�؉�?�q�q�?�q�q�?      �?      �?      �?                      �?              �?              �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�v}hG        hNhG        hNhBKhDKhEh)h,K ��h.��R�(KK��h^�C              �?�t�bhQhchLC       ���R�hgKhhhkKh)h,K ��h.��R�(KK��hL�C       �t�bK��R�}�(hKhuM1hvh)h,K ��h.��R�(KM1��h}�B@L         �                    �?U�ք�?�           ��@              !                   �\@T��_�v�?�            Pw@                                   �?�+$�jP�?$             K@                                 @e@��R[s�?            �A@              
                    �?     ��?             @@                                   X@      �?             @        ������������������������       �                     �?               	                    �M@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?                                  �S@؇���X�?             <@                                   �?      �?	             0@       ������������������������       �                     (@                                  @]@      �?             @        ������������������������       �                     �?        ������������������������       �                     @                                ����?      �?	             (@                                 `\@"pc�
�?             &@                                 @Z@�����H�?             "@                                 �[@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @                                   �J@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @                                  @V@�}�+r��?             3@       ������������������������       �                     $@                                   i@�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        "       #                 ���ٿ�Z�0���?�            �s@        ������������������������       �                      @        $       -                    I@F�F��?�            �s@        %       (                     J@��+7��?             7@       &       '                 �����@4և���?             ,@        ������������������������       �                     �?        ������������������������       �        
             *@        )       *                    �K@X�<ݚ�?             "@        ������������������������       �                     @        +       ,                   �]@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        .       �                   pq@��k�Or�?�            `r@       /       H                   �]@L6�E�i�?�            �l@        0       1                   �`@"Ae���?            �G@        ������������������������       �                     @        2       G                 ����?^����?            �E@       3       4                   �Z@���|���?            �@@        ������������������������       �                     @        5       8                   @[@X�<ݚ�?             ;@        6       7                   �c@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        9       >                    @F@�û��|�?             7@        :       ;                   �i@�q�q�?             "@        ������������������������       �                     @        <       =                   �b@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ?       @                   @b@d}h���?             ,@        ������������������������       �                     @        A       B                   Pc@      �?              @        ������������������������       �                      @        C       D                    �G@r�q��?             @        ������������������������       �                      @        E       F                    \@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     $@        I       x                   �?J� ��w�?{             g@       J       c                    @L@��V���?i            �c@       K       b                    �?\#r��?T            �^@       L       M                   �`@�q��/��?E            �X@       ������������������������       �        '             I@        N       Q                   �c@      �?             H@        O       P                   �c@և���X�?             @       ������������������������       �                     @        ������������������������       �                     @        R       ]                   xp@� ��1�?            �D@       S       T                   0e@��a�n`�?             ?@       ������������������������       �                     1@        U       V                    �C@d}h���?
             ,@        ������������������������       �                     @        W       X                   `e@�z�G��?             $@        ������������������������       �                      @        Y       Z                   @b@      �?              @       ������������������������       �                     @        [       \                   �c@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ^       a                   �p@      �?             $@        _       `                    @E@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     8@        d       k                   `j@����X�?            �A@        e       f                   0a@؇���X�?	             ,@        ������������������������       �                     @        g       j                   @f@����X�?             @        h       i                   �e@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        l       s                   Po@�ՙ/�?             5@        m       n                    �M@�q�q�?             "@        ������������������������       �                     @        o       p                    n@      �?             @        ������������������������       �                      @        q       r                    �O@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        t       w                 ����?r�q��?             (@       u       v                   �`@�<ݚ�?             "@        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        y       �                    �?l��
I��?             ;@       z       {                   �a@"pc�
�?             6@        ������������������������       �                     &@        |       }                   �a@���|���?
             &@        ������������������������       �                     �?        ~       �                   0a@�z�G��?	             $@              �                   �l@      �?              @        �       �                   l@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                    @K@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?p�EG/��?(            �O@        �       �                   �r@��Q��?             4@        �       �                    �?�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?        �       �                   �b@�q�q�?             "@        ������������������������       �                     �?        �       �                    b@      �?              @       ������������������������       �                     @        ������������������������       �                      @        �       �                   w@^����?            �E@       �       �                   �\@>A�F<�?             C@        ������������������������       �                      @        �       �                   �r@4?,R��?             B@        �       �                    �?���|���?	             &@       �       �                    b@      �?              @        �       �                   @`@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                   �b@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �b@`2U0*��?             9@        ������������������������       �                     (@        �       �                   �c@$�q-�?             *@        �       �                   �t@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                     @        �                           �?Nn(����?�            �v@       �       �                   `o@��/���?�            p@       �       �                    @4jf�S�?b            �d@       �       �                 033�?X�n�?P            �`@       �       �                   �e@$�ݏ^��?9            �V@       �       �                   P`@PN���?8            @V@       �       �                   �^@(2��R�?%            �M@       �       �                 033�?P���Q�?             D@       ������������������������       �                     :@        �       �                   �[@؇���X�?             ,@        ������������������������       �                     "@        �       �                   `]@���Q��?             @        ������������������������       �                     �?        �       �                    I@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   P`@�����?             3@        �       �                 ����?X�<ݚ�?             "@       �       �                   @j@����X�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        �       �                   �h@ףp=
�?             $@        �       �                   `@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �m@�q�q�?             >@       �       �                   �i@���Q��?             9@        �       �                 033�?z�G�z�?             $@        �       �                   `h@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                   k@��S���?	             .@        ������������������������       �                     @        �       �                    �G@���|���?             &@        ������������������������       �                     @        �       �                   �a@և���X�?             @        ������������������������       �                      @        �       �                   �m@z�G�z�?             @        ������������������������       �                     @        �       �                   @_@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                    b@�&!��?            �E@       �       �                    �?�q�q�?            �C@        �       �                 033�?      �?              @       �       �                    i@      �?             @        ������������������������       �                      @        �       �                   �a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                   @n@r֛w���?             ?@       �       �                 `ff�?V�a�� �?             =@        ������������������������       �                     @        �       �                    �?�θ�?             :@       �       �                   �_@"pc�
�?
             6@       �       �                   �_@����X�?             ,@        ������������������������       �                      @        �       �                    �I@r�q��?             (@        �       �                   �\@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                      @        �       �                   @`@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                    o@<���D�?            �@@       �       �                   �b@     ��?             @@       �       �                    �? ��WV�?             :@        �       �                    \@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     6@        �       �                   `c@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �                          �?@S�)�q�?7            �V@        �                         `c@�t����?             1@       �                         h~@z�G�z�?             .@       �                          @`@$�q-�?             *@        ������������������������       �                     @                                8s@؇���X�?             @       ������������������������       �                     @                                hv@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @                              ����?�MI8d�?)            �R@        	                          K@�ՙ/�?             5@        
                        �s@ףp=
�?             $@       ������������������������       �                     @                                 �I@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                0b@���|���?             &@                                �L@      �?              @        ������������������������       �                     @                                 a@z�G�z�?             @                                xs@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @                                �`@�NW���?            �J@                                 �?������?             1@                               Pe@$�q-�?	             *@       ������������������������       �                     (@        ������������������������       �                     �?                                �b@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     B@        !      0                   �R@�q-�??             Z@       "      +                ����?p�eU}�?>            �Y@        #      *                  `c@�>4և��?             <@       $      )                  �c@�E��ӭ�?
             2@       %      &                   n@������?	             1@       ������������������������       �                     &@        '      (                  �z@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     $@        ,      -                   @O@�}��L�?.            �R@       ������������������������       �                    �E@        .      /                   @      �?             @@       ������������������������       �                     ?@        ������������������������       �                     �?        ������������������������       �                     �?        �t�bh�h)h,K ��h.��R�(KM1KK��h^�B  ᓔ��?�5�;��?�q����?$�����?B{	�%��?/�����?PuPu�?X|�W|��?      �?      �?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?�$I�$I�?۶m۶m�?      �?      �?              �?      �?      �?      �?                      �?      �?      �?F]t�E�?/�袋.�?�q�q�?�q�q�?�������?�������?      �?                      �?              �?      �?      �?      �?                      �?      �?              �?        (�����?�5��P�?              �?�q�q�?�q�q�?      �?                      �?����?����q�?              �?0�O��?��`=��?Y�B��?zӛ����?�$I�$I�?n۶m۶�?      �?                      �?r�q��?�q�q�?      �?        �������?�������?      �?                      �?���E�?�7�L\��?ł�P���?��e�:}�?�w6�;�?W�+���?              �?�qG��?w�qG��?]t�E]�?F]t�E�?      �?        r�q��?�q�q�?      �?      �?              �?      �?        8��Moz�?��,d!�?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?        I�$I�$�?۶m۶m�?      �?              �?      �?              �?�������?UUUUUU�?      �?              �?      �?      �?                      �?      �?        -d!Y��?Nozӛ��?����?������?��:��?XG��).�?/����?և���X�?      �?              �?      �?۶m۶m�?�$I�$I�?      �?                      �?������?������?�s�9��?�c�1Ƹ?      �?        I�$I�$�?۶m۶m�?      �?        ffffff�?333333�?              �?      �?      �?      �?              �?      �?              �?      �?              �?      �?UUUUUU�?�������?      �?                      �?      �?              �?        �m۶m��?�$I�$I�?۶m۶m�?�$I�$I�?      �?        �m۶m��?�$I�$I�?UUUUUU�?UUUUUU�?      �?                      �?      �?        �<��<��?�a�a�?UUUUUU�?UUUUUU�?              �?      �?      �?      �?              �?      �?      �?                      �?�������?UUUUUU�?9��8���?�q�q�?              �?      �?              �?        Lh/����?h/�����?/�袋.�?F]t�E�?      �?        ]t�E]�?F]t�E�?              �?ffffff�?333333�?      �?      �?      �?      �?      �?                      �?      �?                      �?�������?�������?      �?                      �?�4M�4M�?Y�eY�e�?ffffff�?�������?F]t�E�?]t�E�?              �?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?�qG��?w�qG��?������?Cy�5��?              �?�8��8��?r�q��?]t�E]�?F]t�E�?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?        UUUUUU�?UUUUUU�?              �?      �?        ���Q��?{�G�z�?      �?        �؉�؉�?;�;��?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?�˹�m�?~�Q���?����?w�v�v��?��7�:��?�=�b��?u�՝Vw�?E,�T��?�I��I��?[�[��?B�P�"�?_��׽��?'u_[�?=�"h8��?�������?ffffff�?              �?�$I�$I�?۶m۶m�?              �?�������?333333�?      �?              �?      �?      �?                      �?^Cy�5�?Q^Cy��?r�q��?�q�q�?�m۶m��?�$I�$I�?      �?                      �?              �?�������?�������?      �?      �?              �?      �?                      �?UUUUUU�?UUUUUU�?333333�?�������?�������?�������?      �?      �?              �?      �?              �?        �������?�?              �?]t�E]�?F]t�E�?      �?        ۶m۶m�?�$I�$I�?      �?        �������?�������?              �?      �?      �?              �?      �?              �?              �?        ֔5eMY�?S֔5eM�?UUUUUU�?UUUUUU�?      �?      �?      �?      �?      �?              �?      �?              �?      �?                      �?���{��?�B!��?��{a�?a���{�?      �?        ى�؉��?�؉�؉�?/�袋.�?F]t�E�?�m۶m��?�$I�$I�?              �?�������?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?              �?      �?      �?                      �?              �?              �?|���?|���?      �?      �?;�;��?O��N���?      �?      �?      �?                      �?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        �~�~��?Z�Z��?�������?�������?�������?�������?;�;��?�؉�؉�?              �?�$I�$I�?۶m۶m�?              �?      �?      �?      �?                      �?      �?              �?        L�Ϻ��?��L���?�a�a�?�<��<��?�������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?]t�E]�?F]t�E�?      �?      �?      �?        �������?�������?      �?      �?              �?      �?                      �?      �?        �x+�R�?萚`���?�?xxxxxx�?;�;��?�؉�؉�?              �?      �?              �?      �?              �?      �?                      �?�;�;�?��؉���?��VCӭ?(�J��"�?�m۶m��?�$I�$I�?r�q��?�q�q�?�?xxxxxx�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?O贁N�?�_,�Œ�?              �?      �?      �?              �?      �?              �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJg}�XhG        hNhG        hNhBKhDKhEh)h,K ��h.��R�(KK��h^�C              �?�t�bhQhchLC       ���R�hgKhhhkKh)h,K ��h.��R�(KK��hL�C       �t�bK��R�}�(hKhuM;hvh)h,K ��h.��R�(KM;��h}�B�N         ~                   P`@0����?�           ��@                                   @I@�<ݚ�?�            �s@                                  @h@������?)             L@                                   �?�㙢�c�?             7@                                   �D@      �?              @        ������������������������       �                     �?                                  @[@և���X�?             @        ������������������������       �                     �?        	                           ^@�q�q�?             @        
                            F@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        	             .@                                   �?�eP*L��?            �@@                                   \@      �?             0@                                  @\@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     *@                                  @_@�IєX�?             1@                                  `]@r�q��?             @                                  @H@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     &@               o                    �?�����=�?�            0p@              T                   �`@      �?s            �f@               ?                   �]@�a7���?9            �U@              0                 @33�?Ȩ�I��?!            �J@                #                    �J@�û��|�?             7@        !       "                     J@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        $       %                    W@��S���?
             .@        ������������������������       �                     @        &       /                   �o@�q�q�?             (@       '       (                   @Z@z�G�z�?             $@        ������������������������       �                     @        )       .                    �?�q�q�?             @       *       +                     L@���Q��?             @        ������������������������       �                      @        ,       -                    ^@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        1       :                   �[@r�q��?             >@       2       3                   �_@ףp=
�?             4@       ������������������������       �                     *@        4       9                   �X@����X�?             @       5       6                    �K@      �?             @        ������������������������       �                     �?        7       8                 ����?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ;       <                    \@�z�G��?             $@        ������������������������       �                     �?        =       >                    @O@�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                      @        @       A                    �I@�'�=z��?            �@@        ������������������������       �                      @        B       O                    `@�g�y��?             ?@       C       D                   �Z@������?             1@        ������������������������       �                      @        E       N                   �p@������?             .@       F       M                   �_@8�Z$���?
             *@       G       L                    @O@����X�?             @       H       I                    @L@r�q��?             @       ������������������������       �                     @        J       K                   �^@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        P       S                   Po@d}h���?             ,@       Q       R                    �?      �?              @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        U       n                   0`@��0{9�?:            �W@       V       c                 ����?Ĝ�oV4�?8            �V@        W       b                   `_@��H�}�?             9@       X       Y                    W@���!pc�?             6@        ������������������������       �                     @        Z       a                 hff�?���Q��?             .@       [       \                   @]@�	j*D�?
             *@        ������������������������       �                     @        ]       `                   �T@ףp=
�?             $@        ^       _                   �]@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        d       e                   �b@Pa�	�?(            �P@       ������������������������       �                     C@        f       g                 ����?@4և���?             <@        ������������������������       �                     *@        h       i                    V@�r����?
             .@        ������������������������       �                     �?        j       m                   @c@@4և���?	             ,@        k       l                   �Y@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     @        p       }                    �?l{��b��?1            �S@       q       z                   (r@�LQ�1	�?             G@       r       s                    �?������?            �D@        ������������������������       �                     @        t       y                   �^@ >�֕�?            �A@        u       x                    Y@      �?             0@        v       w                   @V@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     (@        ������������������������       �                     3@        {       |                     L@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                    �@@               �                   �b@�"�,��?	           0z@        �       �                 pff�?F�|����?w             g@        �       �                   Xq@R���Q�?5             T@       �       �                   @d@     ��?-             P@       �       �                   @E@؇���X�?,            �O@        �       �                 �����      �?             @        ������������������������       �                     �?        �       �                   0a@�q�q�?             @        ������������������������       �                     �?        �       �                 ����?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   pa@�^����?(            �M@        ������������������������       �                     2@        �       �                   �j@��r._�?            �D@       �       �                   �^@�d�����?             3@        �       �                     F@և���X�?             @        ������������������������       �                      @        �       �                    �J@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                    �L@r�q��?	             (@       ������������������������       �                     @        �       �                    �?�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                 ����?�C��2(�?             6@       �       �                    �B@�X�<ݺ?             2@        �       �                   �m@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        
             0@        �       �                   �a@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                 @33�?      �?             0@       �       �                   �q@և���X�?             ,@        ������������������������       �                     @        �       �                    �?���Q��?             $@        ������������������������       �                      @        �       �                   @a@      �?              @        ������������������������       �                     �?        �       �                   �`@؇���X�?             @        ������������������������       �                     @        �       �                     J@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                   v@8	C)��?B            @Z@       �       �                   �_@t�F�}�?A            �Y@        �       �                    �?�P�*�?             ?@       �       �                    �D@|��?���?             ;@        ������������������������       �                     @        �       �                 ����?r�q��?             8@        ������������������������       �                     @        �       �                   �j@b�2�tk�?             2@        �       �                    \@����X�?             @        ������������������������       �                      @        �       �                    �I@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                   Pb@"pc�
�?             &@       ������������������������       �                      @        �       �                   �o@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                   p`@@���?T�?+            �Q@        ������������������������       �                     @        �       �                   �j@� y���?*            �P@        �       �                    �?`2U0*��?             9@        ������������������������       �                     *@        �       �                    @J@�8��8��?             (@        �       �                    �I@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     "@        �       �                    @P@���N8�?             E@       �       �                   0a@��G���?            �B@        �       �                    @L@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                   @k@6YE�t�?            �@@        ������������������������       �                     �?        �       �                   �a@      �?             @@       �       �                    @J@������?             .@        �       �                    �?���Q��?             @        ������������������������       �                      @        �       �                   �a@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                 `ff�?ףp=
�?             $@        �       �                    �M@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        
             1@        �       �                    �P@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                   �P@��qM��?�            @m@        �       �                    �?�IєX�?
             1@       ������������������������       �                     *@        �       �                    �?      �?             @        ������������������������       �                      @        �       �                    `@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       :                   @pW�
�?�             k@       �                       833�?r�����?�            �j@       �       �                   �c@�J�ۈ�?S            `a@        �       �                    ]@և���X�?             5@        ������������������������       �                     @        �       �                   `@      �?             0@        �       �                    �?      �?             @        ������������������������       �                     �?        �       �                    @E@���Q��?             @        ������������������������       �                      @        �       �                    @H@�q�q�?             @        ������������������������       �                     �?        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �c@ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        �                         �b@|�9ǣ�?C            �]@                                �n@h�)S;�?=            �[@       ������������������������       �        #            �P@                                 @C@RB)��.�?            �E@                                 �A@���Q��?             @       ������������������������       �                      @        ������������������������       �                     @                                @o@�S����?             C@        ������������������������       �                      @                                s@�����H�?             B@       	                         `@PN��T'�?             ;@       
                         �L@      �?
             0@                                �?؇���X�?             ,@        ������������������������       �                     @                                 �?      �?              @                                @G@����X�?             @        ������������������������       �                     @                                �p@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     &@        ������������������������       �                     "@                                 �?      �?              @        ������������������������       �                     �?                                �c@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @                                Pi@�1��u�?0            @R@        ������������������������       �                     ,@                                �c@L
�q��?*            �M@        ������������������������       �        
             0@               !                   @F@v ��?             �E@        ������������������������       �                     @        "      )                  �c@X�<ݚ�?             B@        #      $                   �H@�����H�?             "@        ������������������������       �                     @        %      (                  �c@z�G�z�?             @       &      '                   �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        *      -                   �H@X�<ݚ�?             ;@        +      ,                hff�?r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        .      /                  �j@�q�q�?             5@        ������������������������       �                      @        0      3                  �p@�d�����?             3@       1      2                   @O@�C��2(�?
             &@       ������������������������       �        	             $@        ������������������������       �                     �?        4      9                   b@      �?              @       5      6                   �K@�q�q�?             @        ������������������������       �                     �?        7      8                   �P@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KM;KK��h^�B�  ���^L�?���Y�?�q�q�?9��8���?n۶m۶�?I�$I�$�?d!Y�B�?�7��Mo�?      �?      �?      �?        ۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?]t�E�?t�E]t�?      �?      �?UUUUUU�?UUUUUU�?              �?      �?              �?        �?�?UUUUUU�?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?F�y�b4�?.�!J��?      �?      �?�qG��?qG�w�?�	�[���?+�R��?��,d!�?8��Moz�?      �?      �?      �?                      �?�?�������?              �?UUUUUU�?UUUUUU�?�������?�������?      �?        UUUUUU�?UUUUUU�?333333�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?                      �?UUUUUU�?�������?�������?�������?              �?�$I�$I�?�m۶m��?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?333333�?ffffff�?      �?        �q�q�?9��8���?              �?      �?        |��|�?|���?      �?        ��{���?�B!��?�?xxxxxx�?              �?�?wwwwww�?;�;��?;�;��?�$I�$I�?�m۶m��?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?      �?        I�$I�$�?۶m۶m�?      �?      �?      �?                      �?      �?        L� &W�?m�w6�;�?����?�!�!�?
ףp=
�?{�G�z�?t�E]t�?F]t�E�?              �?�������?333333�?;�;��?vb'vb'�?      �?        �������?�������?      �?      �?      �?                      �?              �?      �?              �?        |���?|���?              �?�$I�$I�?n۶m۶�?              �?�?�������?      �?        �$I�$I�?n۶m۶�?�������?�������?              �?      �?                      �?      �?        �&��jq�?${�ґ�?Y�B��?��Moz��?������?p>�cp�?              �?�A�A�?��+��+�?      �?      �?      �?      �?              �?      �?                      �?              �?�������?�������?              �?      �?                      �?��/�P�?9����^�?bw�#�?<����?�������?�������?      �?      �?۶m۶m�?�$I�$I�?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?        u_[4�?W'u_�?      �?        �ڕ�]��?ە�]���?Cy�5��?y�5���?�$I�$I�?۶m۶m�?      �?        �������?333333�?              �?      �?        �������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?                      �?]t�E�?F]t�E�?��8��8�?�q�q�?      �?      �?      �?                      �?      �?              �?      �?              �?      �?                      �?      �?      �?۶m۶m�?�$I�$I�?              �?333333�?�������?              �?      �?      �?              �?۶m۶m�?�$I�$I�?      �?              �?      �?              �?      �?              �?        S.�R.��?�h��h��?�������?777777�?�Zk����?�RJ)���?	�%����?{	�%���?              �?UUUUUU�?UUUUUU�?      �?        9��8���?�8��8��?�m۶m��?�$I�$I�?      �?        333333�?�������?              �?      �?        F]t�E�?/�袋.�?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?Zas �
�?�'�K=�?      �?        ~5&��?z�rv��?{�G�z�?���Q��?              �?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?                      �?��y��y�?�a�a�?v�)�Y7�?#�u�)��?      �?      �?              �?      �?        e�M6�d�?'�l��&�?      �?              �?      �?�?wwwwww�?333333�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?        �������?�������?      �?      �?              �?      �?                      �?              �?333333�?�������?      �?                      �?      �?        �z��z��?�
��
��?�?�?              �?      �?      �?              �?      �?      �?              �?      �?        �te�2]�?�,j5��?Dj��V��?�V�9�&�?9ÂKe�?����j�?�$I�$I�?۶m۶m�?              �?      �?      �?      �?      �?              �?333333�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?�������?�������?      �?                      �?Jݗ�V�?�A�Iݷ?b�־a�?� O	�?      �?        S֔5eM�?���)k��?�������?333333�?      �?                      �?(������?^Cy�5�?              �?�q�q�?�q�q�?&���^B�?h/�����?      �?      �?۶m۶m�?�$I�$I�?      �?              �?      �?�m۶m��?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?                      �?      �?              �?              �?      �?              �?۶m۶m�?�$I�$I�?              �?      �?        �s�Ν;�?�1bĈ�?      �?        ��V'�?�pR���?      �?        G�w��?qG�w��?      �?        �q�q�?r�q��?�q�q�?�q�q�?              �?�������?�������?      �?      �?              �?      �?                      �?r�q��?�q�q�?UUUUUU�?�������?      �?                      �?UUUUUU�?UUUUUU�?              �?Cy�5��?y�5���?]t�E�?F]t�E�?      �?                      �?      �?      �?UUUUUU�?UUUUUU�?      �?        �������?�������?              �?      �?              �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ	�tlhG        hNhG        hNhBKhDKhEh)h,K ��h.��R�(KK��h^�C              �?�t�bhQhchLC       ���R�hgKhhhkKh)h,K ��h.��R�(KK��hL�C       �t�bK��R�}�(hKhuMhvh)h,K ��h.��R�(KM��h}�B@@         �                 ����?�+	G�?�           ��@                                `ffֿ�ɞ`s�?�            �v@        ������������������������       �                     @               u                    �?�z�G��?�            �v@                                 @E@�.
���?�            �r@                                   @N@d}h���?             <@                                  �L@�q�q�?             2@              	                   �_@d}h���?	             ,@       ������������������������       �                     "@        
                           �G@���Q��?             @        ������������������������       �                     �?                                  �W@      �?             @        ������������������������       �                     �?        ������������������������       �                     @                                   �?      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     $@               N                    @L@��0p'��?�            �p@              A                   hq@�r�.kx�?�            @j@                                 @]@�KM�]�?m            `e@                                  `k@��.k���?	             1@        ������������������������       �                     @                                  �[@���!pc�?             &@       ������������������������       �                     @        ������������������������       �                      @               2                    �G@XI�~�?d            @c@              '                   �h@�^;\��?7            @V@               &                    �F@�GN�z�?             6@              !                   �\@R���Q�?             4@                                   Pe@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        "       #                   `a@��S�ۿ?
             .@       ������������������������       �                     *@        $       %                    b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        (       -                   �f@�����?(            �P@       )       ,                   �[@�g�y��?$             O@        *       +                    m@8�Z$���?             *@       ������������������������       �                     &@        ������������������������       �                      @        ������������������������       �                    �H@        .       1                    l@z�G�z�?             @        /       0                   �a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        3       @                 ����?��ɉ�?-            @P@       4       7                   `]@ �q�q�?#             H@        5       6                   `e@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        8       ?                   k@�Ń��̧?             E@        9       :                    _@P���Q�?             4@        ������������������������       �                     $@        ;       >                   �_@ףp=
�?	             $@        <       =                   �a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     6@        ������������������������       �        
             1@        B       C                   �q@�(�Tw��?            �C@        ������������������������       �                     @        D       G                   �]@z�G�z�?            �A@        E       F                    �G@      �?             @       ������������������������       �                      @        ������������������������       �                      @        H       I                    `@�חF�P�?             ?@        ������������������������       �                      @        J       M                   �b@��<b���?
             7@        K       L                   �a@      �?             $@       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     *@        O       t                    @R@�-ῃ�?(            �N@       P       g                   �a@T����1�?'             M@       Q       ^                    �M@��J�fj�?            �B@       R       S                   @Z@p�ݯ��?             3@        ������������������������       �                     @        T       U                   @Z@      �?             0@        ������������������������       �                      @        V       ]                    �?؇���X�?
             ,@       W       X                   �_@r�q��?             (@        ������������������������       �                     @        Y       Z                    `@      �?              @        ������������������������       �                     @        [       \                   �c@���Q��?             @       ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        _       d                   �\@�<ݚ�?             2@        `       a                    �N@      �?             @        ������������������������       �                     �?        b       c                   �`@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        e       f                   @^@؇���X�?             ,@        ������������������������       �                      @        ������������������������       �                     (@        h       o                    �?؇���X�?             5@        i       j                   �c@����X�?             @        ������������������������       �                     @        k       l                   @o@      �?             @        ������������������������       �                     �?        m       n                   Pb@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        p       q                    b@@4և���?             ,@       ������������������������       �                      @        r       s                   �d@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        v       �                   �c@:2vz�M�?#            �N@       w       |                   �_@~���L0�?            �H@        x       {                 ����?$�q-�?             *@       y       z                    @K@ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                     @        }       �                    b@b�2�tk�?             B@       ~       �                 hff�?�eP*L��?             6@              �                   �]@p�ݯ��?
             3@        ������������������������       �                     @        �       �                    a@      �?             0@        �       �                    @F@      �?              @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?؇���X�?	             ,@        �       �                     P@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     &@        �       �                   �`@�8��8��?             (@        ������������������������       �                     @        �       �                   pj@z�G�z�?             @        ������������������������       �                     @        �       �                    @I@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �a@2�K36��?�             w@       �       �                 033�?ά��.��?�            @p@        �       �                   Pi@      �?              @        ������������������������       �                     @        �       �                   �_@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �`@<�T]���?�            �o@       �       �                   �`@������?`            @b@       �       �                    �?������?B            @X@       �       �                   �Q@$��$�L�?6            �S@        ������������������������       �                     �?        �       �                 ����?�:�^���?5            �S@        �       �                    �?���N8�?             5@       �       �                    �?�E��ӭ�?             2@        ������������������������       �                     @        �       �                   @_@X�Cc�?             ,@        ������������������������       �                     @        �       �                     K@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                 pff�?���U�?(            �L@        �       �                 ����?�>����?             ;@       �       �                    �? �q�q�?             8@        �       �                    @K@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     5@        �       �                   �e@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     >@        �       �                   `^@�<ݚ�?             2@        �       �                   @[@      �?              @        ������������������������       �                     @        �       �                   �]@z�G�z�?             @        �       �                   �\@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     $@        �       �                 pff�?@�E�x�?            �H@        �       �                    �Q@�8��8��?             (@       ������������������������       �                     &@        ������������������������       �                     �?        ������������������������       �                    �B@        �       �                   @[@Fmq��?>            �Z@        ������������������������       �                     "@        �       �                    @L@����l�?8            @X@       �       �                 033@�5��?             K@       �       �                    �J@��H�}�?             I@       �       �                   Pm@�G�z��?             D@       �       �                    �F@����X�?             5@        �       �                   �b@      �?              @        ������������������������       �                     @        ������������������������       �                     @        �       �                    @J@8�Z$���?             *@       ������������������������       �                      @        �       �                   �X@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                    �H@�S����?	             3@       ������������������������       �                     *@        �       �                    �I@      �?             @       �       �                    �?���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                     @        �       �                   �`@>��C��?            �E@        ������������������������       �                      @        �       �                   0b@� ��1�?            �D@        ������������������������       �        
             .@        �       �                    @M@�	j*D�?             :@        ������������������������       �                     $@        �       �                    �?      �?             0@       �       �                   xu@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �                           �R@�e/
�?I             [@       �       �                   �b@$	4�}�?H            �Z@        ������������������������       �                     ;@        �       �                    �?R���Q�?4             T@        �       �                 ���@������?             1@       �       �                    V@���|���?             &@        ������������������������       �                     �?        �       �                    @M@�z�G��?             $@        ������������������������       �                      @        �       �                 033@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   Pc@�? Da�?(            �O@        �       �                   pc@����X�?             <@       �       �                   P`@�LQ�1	�?             7@       �       �                   pk@��S�ۿ?
             .@        ������������������������       �                     @        �       �                   �l@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    c@      �?              @       ������������������������       �                     @        �       �                   �`@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                    �A@        ������������������������       �                     �?        �t�b��"     h�h)h,K ��h.��R�(KMKK��h^�B  ��C�l�?z?+^���?mާ�d�?&C��6��?              �?ffffff�?333333�?!�M�/�?~���6@�?۶m۶m�?I�$I�$�?UUUUUU�?UUUUUU�?۶m۶m�?I�$I�$�?              �?333333�?�������?              �?      �?      �?              �?      �?              �?      �?      �?                      �?              �?�&�U��?e��?L��K���?�����?�k(���?(�����?�������?�?      �?        t�E]t�?F]t�E�?      �?                      �?5�wL��?V~B����?ҏ~���?p�\��?�袋.��?]t�E�?333333�?333333�?333333�?�������?              �?      �?        �������?�?      �?              �?      �?              �?      �?                      �?g��1��?���@��?��{���?�B!��?;�;��?;�;��?      �?                      �?      �?        �������?�������?      �?      �?      �?                      �?      �?        ?�?��? �����?�������?UUUUUU�?�������?UUUUUU�?      �?                      �?��<��<�?�a�a�?ffffff�?�������?      �?        �������?�������?      �?      �?              �?      �?              �?              �?              �?        �o��o��?� � �?              �?�������?�������?      �?      �?              �?      �?        �Zk����?��RJ)��?      �?        ��,d!�?��Moz��?      �?      �?              �?      �?              �?        �).�u�?�����?�FX�i��?�rO#,��?�"�u�)�?к����?Cy�5��?^Cy�5�?      �?              �?      �?      �?        �$I�$I�?۶m۶m�?UUUUUU�?�������?              �?      �?      �?              �?�������?333333�?      �?                      �?              �?9��8���?�q�q�?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?۶m۶m�?�$I�$I�?              �?      �?        ۶m۶m�?�$I�$I�?�m۶m��?�$I�$I�?      �?              �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?n۶m۶�?�$I�$I�?      �?        �������?UUUUUU�?              �?      �?                      �?��!XG�?��6�S\�?������?����>4�?;�;��?�؉�؉�?�������?�������?              �?      �?                      �?9��8���?�8��8��?t�E]t�?]t�E�?^Cy�5�?Cy�5��?              �?      �?      �?      �?      �?              �?      �?              �?                      �?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?              �?      �?                      �?UUUUUU�?UUUUUU�?      �?        �������?�������?      �?              �?      �?              �?      �?        ����7��?Y�B���?~�~��?�~�~�?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?�������?AA�?�lٲe˶?iҤI�&�? tT����?|q���
�?�3���?��]-n��?      �?        �o��o��?� � �?��y��y�?�a�a�?r�q��?�q�q�?              �?�m۶m��?%I�$I��?              �?�m۶m��?�$I�$I�?              �?      �?                      �?p�}��?	�#����?h/�����?�Kh/��?UUUUUU�?�������?UUUUUU�?UUUUUU�?      �?                      �?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?�q�q�?9��8���?      �?      �?              �?�������?�������?      �?      �?      �?                      �?      �?                      �?9/���?և���X�?UUUUUU�?UUUUUU�?              �?      �?                      �?~�	�[�?�x+�R�?              �?��Id��?2���$�?h/�����?/�����?{�G�z�?
ףp=
�?�������?�������?�$I�$I�?�m۶m��?      �?      �?              �?      �?        ;�;��?;�;��?              �?�������?333333�?              �?      �?        (������?^Cy�5�?      �?              �?      �?333333�?�������?      �?                      �?              �?      �?                      �?qG�w��?$�;��?      �?        ������?������?              �?;�;��?vb'vb'�?              �?      �?      �?�q�q�?�q�q�?              �?      �?              �?        	�%��о?_B{	�%�?�@�Ե�?��bEi�?              �?333333�?333333�?�?xxxxxx�?F]t�E�?]t�E]�?      �?        333333�?ffffff�?      �?              �?      �?              �?      �?                      �?AA�?�������?�$I�$I�?�m۶m��?Y�B��?��Moz��?�?�������?              �?      �?      �?      �?                      �?      �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�ޡhG        hNhG        hNhBKhDKhEh)h,K ��h.��R�(KK��h^�C              �?�t�bhQhchLC       ���R�hgKhhhkKh)h,K ��h.��R�(KK��hL�C       �t�bK��R�}�(hKhuM9hvh)h,K ��h.��R�(KM9��h}�B@N         v                   �`@6������?�           ��@                                  �f@� o�̞�?�            �s@                                  �Z@0w-!��?E             Y@        ������������������������       �                     9@                                  �Z@�7�QJW�?3            �R@        ������������������������       �                      @                                hff�?v���a�?2            @R@                                   �?     ��?             0@       	                           �?�	j*D�?             *@       
                          ``@      �?              @        ������������������������       �                     @                                  `a@z�G�z�?             @        ������������������������       �                     @                                   b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @                                  P`@l�b�G��?%            �L@                                  �?�����H�?             B@                                   _@      �?
             0@                                  �N@�8��8��?             (@       ������������������������       �                     &@        ������������������������       �                     �?                                   �G@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     4@        ������������������������       �                     5@               _                    �?༉p��?�            �j@              X                 ����?�����?c            `b@               K                    @O@rOP\6�?2            @S@       !       .                    �G@���h%��?(            �O@        "       -                    �?��.k���?
             1@       #       &                    �F@X�Cc�?             ,@        $       %                   �y@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        '       ,                    �?և���X�?             @       (       )                    _@�q�q�?             @        ������������������������       �                     @        *       +                   �l@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        /       @                   Hp@��+7��?             G@       0       1                    �?\-��p�?             =@        ������������������������       �                     @        2       3                    @J@"pc�
�?             6@        ������������������������       �                     "@        4       ?                    �?�	j*D�?	             *@       5       >                    @M@      �?             (@       6       =                    �?և���X�?             @       7       <                    �?�q�q�?             @       8       9                   �h@���Q��?             @        ������������������������       �                      @        :       ;                     L@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        A       D                   �]@��.k���?             1@        B       C                    Y@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        E       F                   @_@�z�G��?             $@        ������������������������       �                      @        G       H                    �K@      �?              @        ������������������������       �                      @        I       J                    `@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        L       S                     Q@X�Cc�?
             ,@       M       N                    �?      �?              @        ������������������������       �                      @        O       P                 ����?r�q��?             @        ������������������������       �                     @        Q       R                    V@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        T       U                 ����?�q�q�?             @        ������������������������       �                     �?        V       W                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        Y       ^                    �R@��?^�k�?1            �Q@       Z       [                    `P@@	tbA@�?0            @Q@       ������������������������       �        *             O@        \       ]                    �P@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        `       m                   �`@��v����?*            �P@        a       b                   @Z@�+e�X�?             9@        ������������������������       �                     @        c       d                    �?�����?             3@        ������������������������       �                     @        e       l                    �?     ��?             0@       f       g                   `\@d}h���?             ,@        ������������������������       �                     �?        h       k                     O@8�Z$���?             *@       i       j                    @M@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        n       o                   `c@@4և���?             E@       ������������������������       �                     8@        p       q                    �I@r�q��?             2@        ������������������������       �                      @        r       u                   �h@      �?	             0@        s       t                   �d@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     *@        w       �                 ����?��y�3��?           @z@       x       �                   �g@���@��?�            0p@       y       �                   @E@
�?�            �o@        z                        ����?�	j*D�?             *@       {       ~                   �a@"pc�
�?             &@        |       }                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        �       �                   @b@"pc�
�?�            @n@        �       �                    �?     ��?*             P@       �       �                    �J@ܷ��?��?%             M@        ������������������������       �                     9@        �       �                   p@"pc�
�?            �@@       �       �                 ����? �Cc}�?             <@       �       �                    �?     ��?
             0@       �       �                   Pa@$�q-�?             *@        ������������������������       �                     @        �       �                    �K@؇���X�?             @        �       �                   �a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �g@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     (@        �       �                    �M@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                   �o@���*~�?p            @f@       �       �                   �c@�ȼB���?J            �[@        �       �                    b@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �f@�u��R�?H            �Z@        �       �                    �?�+e�X�?             9@       �       �                    �I@���Q��?	             .@       �       �                    �?�����H�?             "@        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �f@r�q��?             @       �       �                    @M@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     $@        �       �                 833�?ĴF���?8            �T@       �       �                   �b@��(\���?6             T@       �       �                    �?�kb97�?4            @S@       �       �                   �\@���(-�?1            @R@        �       �                    �G@�θ�?             *@       �       �                   �Z@�z�G��?             $@        ������������������������       �                     @        �       �                   �i@      �?             @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �        &             N@        �       �                   �d@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   �c@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �]@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   `]@��y�:�?&            �P@        �       �                   Pc@      �?	             ,@        ������������������������       �                     @        �       �                    �I@���|���?             &@       �       �                   hp@�q�q�?             @        ������������������������       �                     �?        �       �                   �[@z�G�z�?             @        ������������������������       �                      @        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                 ����?�#ʆA��?            �J@       �       �                    @L@t�F�}�?            �I@       �       �                    `@��s����?             E@       �       �                   �_@�q�q�?             5@       �       �                    �E@      �?	             0@       �       �                     E@���|���?             &@       �       �                   �q@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                   �d@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                   �b@���N8�?
             5@        ������������������������       �                     �?        ������������������������       �        	             4@        �       �                   r@�q�q�?             "@        ������������������������       �                      @        �       �                   pe@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    d@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �                         �b@���ѽ��?k             d@        �                          �?R���Q�?4             T@       �       �                   �U@�q�q�?&             K@        ������������������������       �                      @        �       �                   �`@�	j*D�?%             J@        ������������������������       �                     �?        �       
                  �b@�t����?$            �I@       �                          @L@(���@��?!            �G@       �                          @��S���?             >@       �       �                   @_@�û��|�?             7@        �       �                    �D@�<ݚ�?             "@        ������������������������       �                      @        ������������������������       �                     @        �       �                   �V@      �?             ,@        ������������������������       �                     @        �       �                 ����?���|���?	             &@        �       �                    �?���Q��?             @        ������������������������       �                     �?        �       �                    a@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �a@r�q��?             @        ������������������������       �                     �?        �                         �a@z�G�z�?             @       �       �                    �?      �?             @        ������������������������       �                     �?        �                          @e@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @              	                `ff�?�IєX�?             1@                                 @O@r�q��?             @                                �p@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     &@        ������������������������       �                     @        ������������������������       �                     :@              8                   @|��?���?7            @T@                               c@�Z4���?.            �P@        ������������������������       �                     @                                 \@Nd^����?)            �N@                              ����?r�q��?             @                                �Z@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @              7                  0s@���|���?%            �K@             2                  `q@ڡR����?!            �H@             1                   @P@�z�G��?             D@             "                  �j@�d�����?             C@                                 a@��
ц��?	             *@                                �?r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?                                pi@؇���X�?             @        ������������������������       �                     @               !                  @j@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        #      (                  Pc@�J�4�?             9@        $      '                   b@���Q��?             @       %      &                   �F@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        )      *                   �?P���Q�?             4@        ������������������������       �                     $@        +      0                    J@ףp=
�?             $@        ,      -                  Pd@�q�q�?             @        ������������������������       �                     �?        .      /                  �`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        3      4                  `r@�����H�?             "@       ������������������������       �                     @        5      6                  �r@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        	             ,@        �t�bh�h)h,K ��h.��R�(KM9KK��h^�B�  ��X�5�?��S�$e�?b��x�Y�?��a���?�p=
ף�?ףp=
��?              �?0��b�/�?t�@�t�?      �?        �4iҤI�?ٲe˖-�?      �?      �?;�;��?vb'vb'�?      �?      �?              �?�������?�������?      �?              �?      �?              �?      �?                      �?      �?        p�}��?�Gp��?�q�q�?�q�q�?      �?      �?UUUUUU�?UUUUUU�?              �?      �?              �?      �?              �?      �?                      �?              �?p�_���?H&�;u-�?q�{���?G-B���?��O����?dj`��?v]�u]��?EQEQ�?�������?�?%I�$I��?�m۶m��?۶m۶m�?�$I�$I�?      �?                      �?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?zӛ����?Y�B��?a����?�{a���?      �?        /�袋.�?F]t�E�?      �?        vb'vb'�?;�;��?      �?      �?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?333333�?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?      �?                      �?�������?�?�$I�$I�?�m۶m��?      �?                      �?ffffff�?333333�?      �?              �?      �?              �?�������?UUUUUU�?      �?                      �?�m۶m��?%I�$I��?      �?      �?              �?UUUUUU�?�������?              �?      �?      �?              �?      �?        UUUUUU�?UUUUUU�?              �?�������?�������?      �?                      �?�A�A�?_�_��?ہ�v`��?�%~F��?              �?�$I�$I�?۶m۶m�?      �?                      �?      �?        *g��1�?5&����?���Q��?R���Q�?              �?^Cy�5�?Q^Cy��?      �?              �?      �?۶m۶m�?I�$I�$�?      �?        ;�;��?;�;��?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?�$I�$I�?n۶m۶�?              �?UUUUUU�?�������?      �?              �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?��	��	�?�~��~��?L�Ϻ��?к����?YYYYYY�?�������?;�;��?vb'vb'�?F]t�E�?/�袋.�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        /�袋.�?F]t�E�?      �?      �?��=���?a���{�?      �?        /�袋.�?F]t�E�?%I�$I��?۶m۶m�?      �?      �?�؉�؉�?;�;��?      �?        ۶m۶m�?�$I�$I�?      �?      �?              �?      �?              �?        UUUUUU�?UUUUUU�?      �?                      �?      �?        �������?333333�?              �?      �?              �?        ���d%+�?��MmjS�?3���+c�?5'��Ps�?      �?      �?      �?                      �?�@�Ե�?7��XQ�?R���Q�?���Q��?333333�?�������?�q�q�?�q�q�?              �?      �?        UUUUUU�?�������?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?        E�JԮD�?ە�]�ڵ?�������?333333�?�Y�	qV�?�cj`?��իW��?�P�B�
�?ى�؉��?�؉�؉�?ffffff�?333333�?      �?              �?      �?              �?      �?              �?              �?              �?      �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?              �?      �?      �?                      �?�@��~�?~5&��?      �?      �?              �?]t�E]�?F]t�E�?UUUUUU�?UUUUUU�?      �?        �������?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?        e�Cj���?5�x+��?777777�?�������?z��y���?�a�a�?UUUUUU�?UUUUUU�?      �?      �?]t�E]�?F]t�E�?      �?      �?              �?      �?                      �?      �?        �������?333333�?              �?      �?        ��y��y�?�a�a�?              �?      �?        UUUUUU�?UUUUUU�?      �?        �$I�$I�?۶m۶m�?              �?      �?              �?      �?              �?      �?              �?      �?      �?                      �?�싨���?�	���?�������?�������?UUUUUU�?UUUUUU�?      �?        ;�;��?vb'vb'�?      �?        �������?�������?R�٨�l�?W�+���?�������?�?8��Moz�?��,d!�?9��8���?�q�q�?              �?      �?              �?      �?              �?]t�E]�?F]t�E�?�������?333333�?      �?              �?      �?      �?                      �?�������?UUUUUU�?      �?        �������?�������?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?�?�?UUUUUU�?�������?      �?      �?      �?                      �?              �?              �?              �?              �?{	�%���?	�%����?\�՘H�?IT�n��?      �?        �u�y���?���:�?UUUUUU�?�������?UUUUUU�?UUUUUU�?      �?                      �?              �?]t�E]�?F]t�E�?����S��?����X�?ffffff�?333333�?Cy�5��?y�5���?�;�;�?�؉�؉�?UUUUUU�?�������?              �?      �?        ۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?        �z�G��?{�G�z�?�������?333333�?UUUUUU�?UUUUUU�?              �?      �?                      �?ffffff�?�������?      �?        �������?�������?UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?      �?                      �?�q�q�?�q�q�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJQY%hG        hNhG        hNhBKhDKhEh)h,K ��h.��R�(KK��h^�C              �?�t�bhQhchLC       ���R�hgKhhhkKh)h,K ��h.��R�(KK��hL�C       �t�bK��R�}�(hKhuM3hvh)h,K ��h.��R�(KM3��h}�B�L                            �?�Z���?�           ��@              e                   P`@�N��[��?t           �@                                   �? ��r�T�?�             m@                                  �a@��Sݭg�?            �C@              
                    �P@J�8���?             =@              	                   �k@��2(&�?             6@                                  `j@���!pc�?             &@       ������������������������       �                      @        ������������������������       �                     @        ������������������������       �        	             &@        ������������������������       �                     @        ������������������������       �                     $@               "                   0b@.��Zr��?~            @h@                                   �E@8�Z$���?#             J@        ������������������������       �                     �?                                  �]@L紂P�?"            �I@                                  �?`Jj��?             ?@                               hff�?ףp=
�?             4@                                   J@�<ݚ�?             "@        ������������������������       �                     �?                                ����?      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                     &@                                   п      �?             4@        ������������������������       �                     @               !                   P`@�t����?             1@                                    @K@����X�?             @                                  �^@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     $@        #       T                 pff�?.}Z*�?[            �a@       $       %                    �A@���L��?1            �S@        ������������������������       �                     @        &       C                   l@L�qA��?0            �R@       '       4                   �h@�p ��?            �D@        (       /                   @^@�q�q�?             2@        )       .                     M@      �?              @       *       -                    �?r�q��?             @       +       ,                   @]@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        0       3                   `g@ףp=
�?             $@        1       2                    �G@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        5       6                   �V@�LQ�1	�?             7@        ������������������������       �                      @        7       B                    d@����X�?             5@       8       A                   Pk@���y4F�?
             3@       9       :                    @G@�	j*D�?             *@        ������������������������       �                      @        ;       >                   �j@"pc�
�?             &@       <       =                    `@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        ?       @                   �j@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        D       S                   �t@H�V�e��?             A@       E       P                    �N@��� ��?             ?@       F       O                   �a@@4և���?             <@       G       H                   `^@�C��2(�?             6@       ������������������������       �        
             .@        I       J                 ����?����X�?             @        ������������������������       �                     @        K       L                   @_@�q�q�?             @        ������������������������       �                     �?        M       N                   �`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        Q       R                   �q@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        U       ^                   �_@     ��?*             P@        V       W                   e@     ��?	             0@        ������������������������       �                      @        X       ]                    �?d}h���?             ,@       Y       Z                    �K@�8��8��?             (@       ������������������������       �                     $@        [       \                    \@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        _       `                    `P@ �q�q�?!             H@       ������������������������       �                    �D@        a       b                   Pb@����X�?             @        ������������������������       �                     @        c       d                    @�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        f                       ��� @�3_�4��?�            �u@       g       �                    �?zC�Q8��?�            t@       h       �                   �n@�c�w<h�?�            �q@       i       �                   �a@V�a�� �?b             b@       j       o                    �?�1iJ�?X             `@        k       l                   �f@����X�?
             ,@        ������������������������       �                      @        m       n                   �b@r�q��?             (@        ������������������������       �                      @        ������������������������       �                     $@        p       �                 ����?n�����?N            �\@       q       t                    @A@�Zl�i��?7            @T@        r       s                   �c@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        u       �                    @J@�:�^���?4            �S@       v       }                   �[@H%u��?"             I@        w       x                   �Z@�	j*D�?
             *@        ������������������������       �                     @        y       z                   pb@X�<ݚ�?             "@        ������������������������       �                     @        {       |                   �c@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ~       �                   �f@@-�_ .�?            �B@               �                   �f@�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     <@        �       �                 @33�?h�����?             <@       �       �                   @f@���7�?             6@        �       �                   �e@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     2@        ������������������������       �                     @        �       �                    �J@�t����?             A@       �       �                 ����?>���Rp�?             =@        �       �                   @[@      �?              @        ������������������������       �                      @        �       �                 pff�?�q�q�?             @        ������������������������       �                      @        �       �                   @b@      �?             @        ������������������������       �                     �?        �       �                   @c@�q�q�?             @        ������������������������       �                     �?        �       �                 ����?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 033�?؇���X�?             5@        ������������������������       �                     @        �       �                   �`@@�0�!��?
             1@       �       �                   pi@@4և���?             ,@        �       �                    @I@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                   @b@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?���Q��?             @       �       �                   �j@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                    l@      �?
             0@       �       �                    @I@�<ݚ�?             "@        ������������������������       �                     @        �       �                   �b@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        �       �                   Pc@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �C@�f4���?Q             a@        �       �                   �e@�q�q�?	             (@       �       �                    @@@z�G�z�?             $@        ������������������������       �                     �?        �       �                   @a@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �a@J��	�y�?H            @_@        �       �                   �p@�q�q�?             ;@        �       �                   �o@؇���X�?             ,@        �       �                   0o@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     "@        �       �                    �H@��
ц��?	             *@        �       �                   �`@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                 ����?      �?              @       �       �                   pa@���Q��?             @        ������������������������       �                      @        �       �                   a@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                 ����?d}h���?9            �X@       �       �                    o@��3E��?5            @W@        �       �                     K@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �g@r�q��?3            �V@       �       �                   �a@4\�����?2            @V@       �       �                     R@L������?(            @R@       �       �                   d@���Hx�?'             R@        �       �                   r@�(\����?             D@       ������������������������       �        
             8@        �       �                    ]@      �?	             0@        �       �                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     (@        �       �                   0d@     ��?             @@        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 ����?\-��p�?             =@       �       �                 ����?�>����?             ;@       �       �                   Pe@�8��8��?             8@        ������������������������       �                     &@        �       �                     H@8�Z$���?             *@        ������������������������       �                     @        �       �                   @`@      �?              @       �       �                    �J@�q�q�?             @        ������������������������       �                     �?        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �b@      �?
             0@        ������������������������       �                     @        �       �                    �?�C��2(�?             &@        �       �                 ����?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �c@z�G�z�?             @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       
                   �?$�q-�?            �C@       �       �                   pa@ >�֕�?            �A@        ������������������������       �                     $@        �       �                   �\@HP�s��?             9@        ������������������������       �                     @                                  T@ףp=
�?             4@                                 d@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @              	                  `^@�IєX�?
             1@                                0l@r�q��?             @        ������������������������       �                      @                                �c@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     &@                                 �K@      �?             @       ������������������������       �                     @        ������������������������       �                     �?                                �Z@H%u��?             9@        ������������������������       �                      @                                �f@�nkK�?             7@       ������������������������       �                     6@        ������������������������       �                     �?                              ����?��ѝ-�?g            `c@                                �i@�q����?"            �J@       ������������������������       �                     <@                              ����?��H�}�?             9@                               �b@8�A�0��?             6@                               p@�����?             3@        ������������������������       �                     $@                                �p@�q�q�?             "@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @              2                   �R@�IєX�?E            �Y@              '                   �?��^M}�?D            @Y@        !      &                  �c@�<ݚ�?             "@       "      %                   b@���Q��?             @       #      $                   @K@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        (      -                `ff@hl �&�?=             W@       )      *                   �L@����ȫ�?7            �T@        ������������������������       �                     D@        +      ,                  0x@�Ń��̧?             E@       ������������������������       �                    �D@        ������������������������       �                     �?        .      /                   @O@z�G�z�?             $@       ������������������������       �                     @        0      1                   b@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     �?        �t�bh�h)h,K ��h.��R�(KM3KK��h^�B0  �H���x�?����C�?����v�?xP� �?�6�����?����?�i�i�?�|˷|��?|a���?�rO#,��?t�E]t�?��.���?t�E]t�?F]t�E�?              �?      �?                      �?      �?                      �?T���t�?�:*���?;�;��?;�;��?      �?        �������?�������?�B!��?���{��?�������?�������?�q�q�?9��8���?      �?              �?      �?              �?      �?                      �?              �?      �?      �?      �?        �?<<<<<<�?�$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?�
��V�?�z2~���?�4H�4H�?��o��o�?              �?t�@��?�K~���?8��18�?dp>�c�?UUUUUU�?UUUUUU�?      �?      �?UUUUUU�?�������?      �?      �?      �?                      �?              �?      �?        �������?�������?UUUUUU�?UUUUUU�?              �?      �?              �?        d!Y�B�?Nozӛ��?      �?        �$I�$I�?�m۶m��?(������?6��P^C�?;�;��?vb'vb'�?      �?        F]t�E�?/�袋.�?�q�q�?�q�q�?              �?      �?              �?      �?      �?                      �?              �?      �?        iiiiii�?ZZZZZZ�?�{����?�B!��?n۶m۶�?�$I�$I�?]t�E�?F]t�E�?      �?        �m۶m��?�$I�$I�?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?      �?     ��?      �?      �?      �?        ۶m۶m�?I�$I�$�?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?              �?        UUUUUU�?�������?              �?�$I�$I�?�m۶m��?              �?UUUUUU�?UUUUUU�?      �?                      �?�avp��?�<���?�c�Ka�??q��z��?��c-C�?ƟH8�y�?��{a�?a���{�?���+��?uE]QW��?�m۶m��?�$I�$I�?              �?�������?UUUUUU�?              �?      �?        �K*���?A�V���?�"e����?�����H�?UUUUUU�?UUUUUU�?              �?      �?        � � �?�o��o��?)\���(�?���Q��?vb'vb'�?;�;��?      �?        r�q��?�q�q�?      �?        �������?�������?              �?      �?        S�n0E�?к����?9��8���?�q�q�?      �?                      �?      �?        �m۶m��?�$I�$I�?�.�袋�?F]t�E�?      �?      �?      �?                      �?      �?              �?        �������?�������?�i��F�?GX�i���?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?۶m۶m�?�$I�$I�?      �?        ZZZZZZ�?�������?n۶m۶�?�$I�$I�?۶m۶m�?�$I�$I�?              �?      �?              �?        UUUUUU�?UUUUUU�?      �?                      �?�������?333333�?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?      �?�q�q�?9��8���?              �?�������?333333�?              �?      �?        ۶m۶m�?�$I�$I�?              �?      �?        ��J��?΂j����?UUUUUU�?UUUUUU�?�������?�������?      �?        �q�q�?�q�q�?              �?      �?              �?        j�t��?+�����?UUUUUU�?UUUUUU�?�$I�$I�?۶m۶m�?�������?333333�?              �?      �?                      �?�;�;�?�؉�؉�?�������?�������?              �?      �?              �?      �?333333�?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?I�$I�$�?۶m۶m�?'�h��&�?f�]v�e�?UUUUUU�?UUUUUU�?      �?                      �?�������?UUUUUU�?�{��^��?B�P�"�?�Ǐ?~�?����?9��8���?9��8��?333333�?�������?      �?              �?      �?      �?      �?              �?      �?              �?              �?      �?UUUUUU�?UUUUUU�?      �?                      �?a����?�{a���?�Kh/��?h/�����?UUUUUU�?UUUUUU�?      �?        ;�;��?;�;��?      �?              �?      �?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?              �?              �?                      �?              �?      �?      �?              �?]t�E�?F]t�E�?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?�������?�������?      �?      �?              �?      �?                      �?�؉�؉�?;�;��?��+��+�?�A�A�?      �?        q=
ףp�?{�G�z�?      �?        �������?�������?UUUUUU�?UUUUUU�?              �?      �?        �?�?�������?UUUUUU�?      �?              �?      �?              �?      �?              �?              �?      �?      �?                      �?���Q��?)\���(�?      �?        d!Y�B�?�Mozӛ�?              �?      �?        +�"�*�?u;T�Cu�?�x+�R�?�Cj��V�?              �?{�G�z�?
ףp=
�?颋.���?/�袋.�?Q^Cy��?^Cy�5�?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        �?�?z��~�X�?�F�tj�?�q�q�?9��8���?�������?333333�?      �?      �?      �?                      �?      �?                      �?Y�B��?ozӛ���?������?������?              �?�a�a�?��<��<�?              �?      �?        �������?�������?              �?      �?      �?              �?      �?              �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ��fbhG        hNhG        hNhBKhDKhEh)h,K ��h.��R�(KK��h^�C              �?�t�bhQhchLC       ���R�hgKhhhkKh)h,K ��h.��R�(KK��hL�C       �t�bK��R�}�(hKhuM5hvh)h,K ��h.��R�(KM5��h}�B@M         �                 ����?�#i����?�           ��@               �                    �? �&�T�?�             w@              �                     R@b��t��?�            �s@              �                 ����? ������?�            @s@              $                    �?��B�?�            �q@                                  �q@�D��?            �H@                                  �J@:�&���?            �C@                                  i@ףp=
�?             4@        	       
                    @A@�q�q�?             @        ������������������������       �                     @                                  pd@�q�q�?             @        ������������������������       �                     �?                                    H@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     ,@                                   @K@�d�����?             3@        ������������������������       �                      @                                  �c@@�0�!��?             1@                                 @_@      �?             0@                                   �N@      �?              @        ������������������������       �                     @                                   k@�q�q�?             @        ������������������������       �                     �?                                  �m@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?                                  �c@���Q��?             $@        ������������������������       �                     @                !                   �_@և���X�?             @        ������������������������       �                      @        "       #                 ����?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        %       6                   `\@�P��G7�?�            @m@        &       5                    �O@�LQ�1	�?             7@       '       4                   �[@����X�?             5@       (       -                   �X@�q�q�?             2@       )       *                   @\@"pc�
�?             &@        ������������������������       �                     �?        +       ,                    �?ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        .       /                   �\@և���X�?             @        ������������������������       �                     �?        0       3                    �M@�q�q�?             @       1       2                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        7       t                   �d@�$
��
�?}            `j@       8       s                   �d@�Zű���?^             d@       9       ^                     L@">R��?]            �c@       :       ]                   pb@�8'��?F            @^@       ;       H                   `g@�����??            �Z@        <       C                   `^@ҳ�wY;�?             1@        =       B                    @J@����X�?             @       >       A                   �e@r�q��?             @        ?       @                   �\@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        D       E                    �J@ףp=
�?             $@       ������������������������       �                      @        F       G                    @K@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        I       \                   �a@ą%�E�?2            @V@       J       [                    �?����?1            �U@       K       T                   �a@ wVX(6�?-            @T@        L       Q                    �J@���B���?             :@       M       N                   0a@P���Q�?             4@       ������������������������       �        	             1@        O       P                    �I@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        R       S                   �^@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        U       Z                    c@h㱪��?            �K@        V       W                   �m@�>����?             ;@       ������������������������       �        	             2@        X       Y                   �[@�<ݚ�?             "@        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     <@        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     .@        _       p                    �N@�d�����?             C@       `       m                    b@և���X�?             5@       a       h                   �`@�q�q�?	             .@       b       c                   �k@X�<ݚ�?             "@        ������������������������       �                      @        d       g                   �_@����X�?             @       e       f                   r@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        i       l                 @33�?r�q��?             @        j       k                   @f@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        n       o                   P`@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        q       r                   @t@�IєX�?             1@       ������������������������       �        
             0@        ������������������������       �                     �?        ������������������������       �                      @        u       |                   pf@HP�s��?             I@       v       w                   q@�7��?            �C@       ������������������������       �                     :@        x       {                   `e@8�Z$���?             *@       y       z                   r@�<ݚ�?             "@        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        }       ~                   �c@"pc�
�?	             &@        ������������������������       �                     �?               �                    @C@ףp=
�?             $@        ������������������������       �                     @        �       �                    @D@z�G�z�?             @        �       �                   @b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �Q@`�Q��?             9@        ������������������������       �                     @        �       �                   �c@�KM�]�?             3@        ������������������������       �                     $@        �       �                   @[@�<ݚ�?             "@        ������������������������       �                     @        �       �                    �?�q�q�?             @       �       �                    @G@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                   �O@~h����?'             L@        ������������������������       �                     6@        �       �                   �p@H�V�e��?             A@       �       �                   �`@ �o_��?             9@        �       �                   @^@r�q��?             @        �       �                   @\@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?�KM�]�?             3@        �       �                    `@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �`@�IєX�?             1@       ������������������������       �                     $@        �       �                 ����?؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        �       �                    �?�������?�            �v@        �       �                   �h@�q�q�?2             R@        �       �                 ����?      �?             4@       �       �                    �L@�θ�?             *@        ������������������������       �                      @        �       �                   �[@���Q��?             @        ������������������������       �                      @        �       �                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �]@ s�n_Y�?%             J@        �       �                   `m@r�q��?             @        �       �                 033@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �K@�LQ�1	�?              G@        �       �                 pff�?      �?              @       �       �                   �a@���Q��?             @        ������������������������       �                      @        �       �                     J@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   0c@�˹�m��?             C@       �       �                    _@h�����?             <@        �       �                    �P@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     5@        �       �                    �?z�G�z�?             $@       �       �                   xu@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        �                       033�?f,��B��?�            `r@       �                         �c@��O5���?u            �h@       �       �                   �\@6�\�{��?g            `e@        �       �                   �X@���N8�?             E@        �       �                   �`@r�q��?             (@       �       �                   �k@�q�q�?             @        ������������������������       �                     �?        �       �                    �K@z�G�z�?             @        ������������������������       �                     @        �       �                   q@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     >@        �                         �e@L�mN�?J             `@       �                         c@�q�q�?G             ^@       �       �                   P`@v�XԖ�?B            �Z@        �       �                    `@�2�o�U�?            �K@       �       �                   @Z@���N8�?             E@        ������������������������       �                     @        �       �                   �R@�E��ӭ�?             B@        �       �                    �N@�X�<ݺ?	             2@       ������������������������       �                     .@        �       �                   �`@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 ����?      �?
             2@       �       �                   �b@���Q��?	             .@       �       �                    �?�	j*D�?             *@       �       �                   `a@      �?             (@       �       �                   �\@և���X�?             @        �       �                    �I@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                    o@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                    �K@��
ц��?             *@        �       �                    �?؇���X�?             @        ������������������������       �                     @        �       �                   �]@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       
                   �R@>a�����?#            �I@       �                       ����?�q��/��?"            �H@        �                          �?�<ݚ�?             2@       �       �                    �?���Q��?	             $@       �       �                    @H@����X�?             @        ������������������������       �                      @        ������������������������       �                     @                                 `X@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @              	                  0b@`Jj��?             ?@                                �?(;L]n�?             >@                                �Q@$�q-�?	             *@        ������������������������       �                     �?        ������������������������       �                     (@        ������������������������       �                     1@        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     ,@                                 @L@X�<ݚ�?             "@        ������������������������       �                     @                                 �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @                                �[@���Q��?             9@        ������������������������       �                     @                              ����?���y4F�?             3@        ������������������������       �                     $@                              033�?X�<ݚ�?             "@        ������������������������       �                      @                                �_@����X�?             @                                �^@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @              0                ��� @@4և���?G            �X@              /                  �c@�LQ�1	�?#             G@             *                   �?Du9iH��?             �E@              )                   �? 	��p�?             =@       !      &                   �M@���}<S�?             7@       "      %                  �X@P���Q�?             4@        #      $                  �`@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �        
             0@        '      (                   �N@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        +      .                   _@@4և���?             ,@        ,      -                  �a@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                     @        1      2                   @O@ pƵHP�?$             J@       ������������������������       �                     F@        3      4                   a@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        �t�b��     h�h)h,K ��h.��R�(KM5KK��h^�BP  �5�;���?%e��?��7��M�?���,d�?}˷|˷�?� � �?�'�Y�	�?j`���?�'�� T�?�`�}��?������??4և���?�A�A�?�o��o��?�������?�������?UUUUUU�?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?              �?        Cy�5��?y�5���?              �?ZZZZZZ�?�������?      �?      �?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?      �?                      �?      �?                      �?�������?333333�?              �?�$I�$I�?۶m۶m�?              �?�������?�������?      �?                      �?Z��Y���?��)��)�?d!Y�B�?Nozӛ��?�$I�$I�?�m۶m��?UUUUUU�?UUUUUU�?F]t�E�?/�袋.�?      �?        �������?�������?              �?      �?        �$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?�������?�������?      �?                      �?              �?              �?      �?        =:�oL�??�A��?Q��/��?��J1Aw�?�X����?ɝ��3 �?N�zv�?�eP*L��?��!5�x�?5�x+��?�������?�������?�$I�$I�?�m۶m��?UUUUUU�?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        �������?�������?      �?              �?      �?              �?      �?        �as���?��g<�?��֡�l�?/�I���?k~X�<�?�<ݚ�?��؉���?ى�؉��?ffffff�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?        UUUUUU�?UUUUUU�?      �?                      �?־a���?��)A��?�Kh/��?h/�����?      �?        9��8���?�q�q�?              �?      �?              �?              �?                      �?      �?        Cy�5��?y�5���?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?r�q��?�q�q�?              �?�m۶m��?�$I�$I�?      �?      �?              �?      �?              �?        �������?UUUUUU�?      �?      �?              �?      �?              �?        UUUUUU�?UUUUUU�?      �?                      �?�?�?      �?                      �?              �?q=
ףp�?{�G�z�?��[��[�?�A�A�?      �?        ;�;��?;�;��?9��8���?�q�q�?              �?      �?              �?        /�袋.�?F]t�E�?              �?�������?�������?      �?        �������?�������?      �?      �?      �?                      �?      �?        ��(\���?{�G�z�?              �?�k(���?(�����?      �?        9��8���?�q�q�?      �?        UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?�m۶m��?%I�$I��?              �?iiiiii�?ZZZZZZ�?
ףp=
�?�Q����?UUUUUU�?�������?      �?      �?              �?      �?                      �?�k(���?(�����?      �?      �?      �?                      �?�?�?      �?        ۶m۶m�?�$I�$I�?              �?      �?              �?        p��Z9��?�D����?�������?�������?      �?      �?ى�؉��?�؉�؉�?      �?        �������?333333�?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?;�;��?�;�;�?�������?UUUUUU�?      �?      �?      �?                      �?      �?        Y�B��?��Moz��?      �?      �?333333�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?                      �?^Cy�5�?��P^Cy�?�$I�$I�?�m۶m��?�$I�$I�?۶m۶m�?              �?      �?                      �?�������?�������?�q�q�?�q�q�?              �?      �?              �?        ŕ�(�?�Z��5;�?��S�r
�?�Cc}�?Fs�e4�?.����2�?�a�a�?��y��y�?UUUUUU�?�������?UUUUUU�?UUUUUU�?      �?        �������?�������?              �?      �?      �?              �?      �?                      �?              �?2g�s��?4�9c��?�������?UUUUUU�?��sHM0�?���s�?�S�<%��?־a��?��y��y�?�a�a�?              �?r�q��?�q�q�?�q�q�?��8��8�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?�������?333333�?;�;��?vb'vb'�?      �?      �?۶m۶m�?�$I�$I�?      �?      �?              �?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?      �?              �?              �?        �;�;�?�؉�؉�?�$I�$I�?۶m۶m�?              �?UUUUUU�?UUUUUU�?              �?      �?              �?        �?�������?և���X�?/����?�q�q�?9��8���?�������?333333�?�$I�$I�?�m۶m��?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?                      �?�B!��?���{��?�?�������?;�;��?�؉�؉�?      �?                      �?              �?      �?              �?                      �?�q�q�?r�q��?              �?�������?�������?              �?      �?        333333�?�������?              �?6��P^C�?(������?      �?        r�q��?�q�q�?              �?�m۶m��?�$I�$I�?UUUUUU�?UUUUUU�?      �?                      �?      �?        �$I�$I�?n۶m۶�?Y�B��?��Moz��?w�qGܱ?qG�w��?�{a���?������?d!Y�B�?ӛ���7�?�������?ffffff�?      �?      �?              �?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?              �?�$I�$I�?n۶m۶�?      �?      �?              �?      �?                      �?      �?        ;�;��?'vb'vb�?              �?      �?      �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ$�phG        hNhG        hNhBKhDKhEh)h,K ��h.��R�(KK��h^�C              �?�t�bhQhchLC       ���R�hgKhhhkKh)h,K ��h.��R�(KK��hL�C       �t�bK��R�}�(hKhuM;hvh)h,K ��h.��R�(KM;��h}�B�N         *                   �_@"��G,�?�           ��@               #                    �?��˥W1�?V            `a@                                   `@��.��?%            �N@                                  `]@`2U0*��?             9@        ������������������������       �                     .@                                   �?ףp=
�?             $@                                  I@؇���X�?             @                                  @N@r�q��?             @       	       
                    �?�q�q�?             @        ������������������������       �                     �?                                  `^@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @                                033�?      �?             B@                                  I@�LQ�1	�?             7@                                  �?����X�?             5@        ������������������������       �                     @                                  �Z@�q�q�?             2@        ������������������������       �                     @                                  �`@�eP*L��?             &@                               ����?      �?              @                                  �]@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @               "                   �\@$�q-�?
             *@                !                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     $@        $       %                    @O@ ���J��?1            �S@       ������������������������       �        (            �L@        &       )                   �`@�����?	             5@        '       (                   `c@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     ,@        +       �                    �I@@�����?h           ��@        ,       �                 033�?L
�q��?�            �m@       -       N                    �E@d,���O�?}            �i@        .       G                   hq@��2(&�?8             V@       /       F                    @D@@4և���?/            �Q@       0       =                    @C@�Ra����?             F@       1       6                   �b@�FVQ&�?            �@@        2       3                   @b@      �?              @        ������������������������       �                     @        4       5                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        7       8                   `f@`2U0*��?             9@       ������������������������       �        
             .@        9       <                   �c@ףp=
�?             $@        :       ;                   �f@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        >       E                   �f@���!pc�?             &@       ?       D                    �C@�����H�?             "@       @       C                   �]@      �?             @        A       B                 @33�?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     :@        H       I                    �?b�2�tk�?	             2@        ������������������������       �                      @        J       K                   �d@     ��?             0@       ������������������������       �                      @        L       M                    �A@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        O       x                   Hq@J�8���?E             ]@       P       w                    @I@���j��?7             W@       Q       r                    �?�w���?0            @T@       R       k                 ����?F�����?+            @R@       S       \                   �]@:ɨ��?&            �P@        T       U                   `Z@�LQ�1	�?             7@        ������������������������       �                     @        V       Y                    �F@      �?	             4@        W       X                   �f@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        Z       [                    �H@$�q-�?             *@       ������������������������       �                     (@        ������������������������       �                     �?        ]       `                   �k@X�EQ]N�?            �E@        ^       _                   �\@���!pc�?             &@        ������������������������       �                     @        ������������������������       �                      @        a       b                 ����?      �?             @@       ������������������������       �                     7@        c       j                   �p@�<ݚ�?             "@       d       i                    b@      �?              @       e       h                 ����?      �?             @       f       g                    �H@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        l       m                   �a@����X�?             @        ������������������������       �                     @        n       o                   @`@�q�q�?             @        ������������������������       �                     �?        p       q                    �G@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        s       t                   @_@      �?              @        ������������������������       �                     @        u       v                    @G@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     &@        y       �                   p`@�q�q�?             8@        z       }                 @33�?����X�?             @        {       |                   �r@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ~                           �?      �?             @        ������������������������       �                     �?        �       �                   `]@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?�t����?	             1@       �       �                   `c@      �?             0@       �       �                   @b@���|���?             &@       �       �                   b@�z�G��?             $@       �       �                    @I@���Q��?             @       ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                   �r@      �?             @@       �       �                   �d@@4և���?             <@        �       �                    �H@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 `ff@`2U0*��?             9@       ������������������������       �                     2@        �       �                   �b@؇���X�?             @        �       �                     H@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �a@      �?             @       ������������������������       �                      @        ������������������������       �                      @        �       $                   �?C nNs�?�            pv@       �                         �a@�\U�a9�?�            r@       �                          @R@��H.��?}             i@       �       �                 ����?$/����?{            `h@        �       �                   �_@���@��?2            �R@        �       �                   @[@��X��?             <@        �       �                   �\@      �?             @        ������������������������       �                      @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                 @33�?      �?             8@       �       �                    e@��s����?             5@       �       �                   `i@R���Q�?             4@        ������������������������       �                     @        ������������������������       �                     1@        ������������������������       �                     �?        �       �                    _@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   pf@*
;&���?             G@        �       �                   @a@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    @L@X�EQ]N�?            �E@        ������������������������       �                     3@        �       �                   �n@�q�q�?             8@        �       �                    _@      �?              @        ������������������������       �                      @        �       �                   �`@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                 ����?      �?	             0@       �       �                   �s@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?2/�o���?I            @^@       �       �                    _@�y�ʍ+�?8             W@        �       �                    �P@$�q-�?             :@       �       �                   �X@ �q�q�?             8@        �       �                    �M@؇���X�?             @        �       �                   �W@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     1@        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �?      �?'            �P@        �       �                 033�?d��0u��?             >@       �       �                    i@�G��l��?             5@        ������������������������       �                      @        �       �                   �a@�\��N��?             3@        ������������������������       �                     @        �       �                   �n@�	j*D�?             *@        ������������������������       �                     @        �       �                    a@X�<ݚ�?             "@       �       �                   h~@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        �       �                 `ff@b�2�tk�?             B@       �       �                   �d@     ��?             @@       �       �                   @_@������?             >@        �       �                 ����?�C��2(�?             &@       �       �                   `k@؇���X�?             @        ������������������������       �                     @        �       �                    �N@      �?             @       �       �                   �o@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    @M@p�ݯ��?             3@       �       �                   �a@��
ц��?             *@       �       �                    �L@�z�G��?             $@       �       �                 ����?և���X�?             @        ������������������������       �                      @        �       �                   �k@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        �       �                    @ܷ��?��?             =@       �       �                   @^@ �q�q�?             8@        �       �                    �?ףp=
�?             $@        �       �                    @L@z�G�z�?             @        ������������������������       �                     @        �       �                   `]@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     ,@                                 p`@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @                                �b@��~l�?0            @V@        ������������������������       �        
             3@                              ����?�z�G��?&            �Q@                                 k@�'�=z��?            �@@        ������������������������       �                     @        	                      ����?և���X�?             <@       
                        �c@�d�����?	             3@                                @m@X�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                     @                                �_@ףp=
�?             $@        ������������������������       �                     @                                a@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @                                �?�<ݚ�?             "@        ������������������������       �                      @                              pff�?����X�?             @        ������������������������       �                     �?                              `ff�?r�q��?             @        ������������������������       �                     @                                pr@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @              #                   �?������?            �B@             "                  0m@r�q��?             8@             !                  l@�	j*D�?             *@                                �c@ףp=
�?             $@       ������������������������       �                     "@        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     &@        ������������������������       �                     *@        %      4                   �P@��R[s�?,            �Q@       &      )                   `@^l��[B�?$             M@        '      (                  hr@�<ݚ�?             "@       ������������������������       �                     @        ������������������������       �                      @        *      +                  ``@�q��/��?            �H@        ������������������������       �                     (@        ,      3                ����?�MI8d�?            �B@        -      2                  �c@      �?
             (@       .      1                   @L@؇���X�?             @        /      0                ����?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     9@        5      :                433�?�q�q�?             (@       6      9                  Pk@      �?              @       7      8                  b@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KM;KK��h^�B�  �UK���?U�)|��?'!����?ۻ��<�?������?�����?{�G�z�?���Q��?              �?�������?�������?�$I�$I�?۶m۶m�?UUUUUU�?�������?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?                      �?              �?              �?      �?      �?d!Y�B�?Nozӛ��?�$I�$I�?�m۶m��?              �?UUUUUU�?UUUUUU�?              �?t�E]t�?]t�E�?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?      �?        ;�;��?�؉�؉�?UUUUUU�?UUUUUU�?      �?                      �?              �?�A�A�?��-��-�?              �?�a�a�?=��<���?�$I�$I�?�m۶m��?              �?      �?                      �? �����?���?��V'�?�pR���?�������?PPPPPP�?��.���?t�E]t�?n۶m۶�?�$I�$I�?]t�E]�?]t�E�?>����?|���?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?���Q��?{�G�z�?      �?        �������?�������?      �?      �?              �?      �?              �?        F]t�E�?t�E]t�?�q�q�?�q�q�?      �?      �?      �?      �?      �?                      �?      �?              �?                      �?      �?        �8��8��?9��8���?      �?              �?      �?      �?              �?      �?      �?                      �?�rO#,��?|a���?ozӛ���?!Y�B�?��Hx��?�n���?�P�B�
�?�^�z���?N6�d�M�?e�M6�d�?d!Y�B�?Nozӛ��?      �?              �?      �?�$I�$I�?۶m۶m�?              �?      �?        ;�;��?�؉�؉�?              �?      �?        w�qG�?qG�wĽ?F]t�E�?t�E]t�?              �?      �?              �?      �?      �?        9��8���?�q�q�?      �?      �?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?                      �?�$I�$I�?�m۶m��?              �?UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?      �?      �?      �?              �?      �?              �?      �?              �?        �������?�������?�m۶m��?�$I�$I�?UUUUUU�?UUUUUU�?              �?      �?              �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?�������?�������?      �?      �?F]t�E�?]t�E]�?333333�?ffffff�?333333�?�������?              �?      �?                      �?      �?                      �?      �?              �?      �?�$I�$I�?n۶m۶�?UUUUUU�?UUUUUU�?      �?                      �?{�G�z�?���Q��?              �?�$I�$I�?۶m۶m�?      �?      �?      �?                      �?              �?      �?      �?              �?      �?        *��M��?k�"Y��?�@�m�?��_�}�?)\���(�?�G�z��? �����?�?�?�?L�Ϻ��?к����?n۶m۶�?%I�$I��?      �?      �?              �?      �?      �?              �?      �?              �?      �?z��y���?�a�a�?333333�?333333�?              �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?        ���,d!�?8��Moz�?UUUUUU�?UUUUUU�?      �?                      �?w�qG�?qG�wĽ?      �?        UUUUUU�?�������?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?              �?      �?      �?      �?      �?                      �?      �?        ��!pc�?�GN��?�,d!Y�?��Moz��?;�;��?�؉�؉�?UUUUUU�?�������?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?      �?      �?              �?      �?              �?      �?wwwwww�?DDDDDD�?1�0��?��y��y�?      �?        �5��P�?y�5���?              �?vb'vb'�?;�;��?      �?        r�q��?�q�q�?�������?�������?              �?      �?              �?                      �?�8��8��?9��8���?      �?      �?wwwwww�?�?]t�E�?F]t�E�?۶m۶m�?�$I�$I�?      �?              �?      �?UUUUUU�?UUUUUU�?              �?      �?              �?              �?        ^Cy�5�?Cy�5��?�؉�؉�?�;�;�?333333�?ffffff�?۶m۶m�?�$I�$I�?      �?        �������?�������?      �?                      �?              �?      �?              �?                      �?              �?a���{�?��=���?UUUUUU�?�������?�������?�������?�������?�������?              �?      �?      �?              �?      �?                      �?              �?�������?333333�?      �?                      �?      �?        ��x�3�?�9�as�?              �?333333�?ffffff�?|��|�?|���?      �?        ۶m۶m�?�$I�$I�?y�5���?Cy�5��?�q�q�?r�q��?              �?      �?        �������?�������?              �?�������?�������?      �?                      �?9��8���?�q�q�?      �?        �m۶m��?�$I�$I�?              �?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?        к����?��g�`��?UUUUUU�?�������?;�;��?vb'vb'�?�������?�������?              �?      �?              �?                      �?              �?PuPu�?X|�W|��?��=���?�=�����?9��8���?�q�q�?      �?                      �?և���X�?/����?              �?L�Ϻ��?��L���?      �?      �?۶m۶m�?�$I�$I�?      �?      �?      �?                      �?      �?                      �?              �?�������?�������?      �?      �?      �?      �?      �?                      �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJW:+LhG        hNhG        hNhBKhDKhEh)h,K ��h.��R�(KK��h^�C              �?�t�bhQhchLC       ���R�hgKhhhkKh)h,K ��h.��R�(KK��hL�C       �t�bK��R�}�(hKhuMhvh)h,K ��h.��R�(KM��h}�B�G         �                    �?�#i����?�           ��@              �                   �a@pٛ'��?r           X�@              p                 033�? � �m$�?           @|@                                 �c@�<ݚ�?�            pq@                                  P`@^������?            �A@                               ����?�S����?             3@                                 @E@�����H�?             2@                                  �?��S�ۿ?             .@       	       
                    `@�C��2(�?	             &@       ������������������������       �                     $@        ������������������������       �                     �?        ������������������������       �                     @                                   �L@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?                                  @_@     ��?	             0@        ������������������������       �                     @                                  `a@�	j*D�?             *@        ������������������������       �                     @                                ����?�q�q�?             @        ������������������������       �                      @                                   b@      �?             @        ������������������������       �                      @        ������������������������       �                      @               Y                 ����?Jy��]0�?�            �n@              :                   �o@�Y{~u4�?w            `h@              '                   �]@|�űN�?L            @]@               &                   �\@      �?             8@                                  �?��<b���?             7@        ������������������������       �                     @                !                    _@ףp=
�?             4@        ������������������������       �                     �?        "       #                   0n@�}�+r��?             3@       ������������������������       �                     1@        $       %                   �[@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        (       -                   �f@����D��?;            @W@        )       *                   �f@P���Q�?             4@       ������������������������       �        
             1@        +       ,                   @_@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        .       /                    `@ �й���?/            @R@        ������������������������       �                     ?@        0       9                   ``@�Ń��̧?             E@       1       2                    �F@���N8�?             5@       ������������������������       �        	             (@        3       8                   0m@�����H�?             "@        4       5                   �Z@�q�q�?             @        ������������������������       �                     �?        6       7                   �j@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     5@        ;       X                    @N@R�}e�.�?+            �S@       <       =                   @[@D˩�m��?)            �R@        ������������������������       �                     �?        >       E                   `]@��oh���?(            @R@        ?       D                   e@��
ц��?             *@       @       C                   Pc@�z�G��?             $@        A       B                     G@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        F       U                    �?r�q��?              N@       G       H                   �^@t�6Z���?            �K@        ������������������������       �        
             0@        I       N                    `@x�����?            �C@        J       M                   �_@      �?              @       K       L                   �d@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        O       P                   �`@��� ��?             ?@        ������������������������       �                     1@        Q       R                   �q@����X�?	             ,@        ������������������������       �                     @        S       T                    �E@      �?              @       ������������������������       �                     @        ������������������������       �                     @        V       W                   Pd@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        Z       o                    @P@�����?            �H@       [       b                    @I@t/*�?            �G@        \       ]                 hff�?�q�q�?             (@        ������������������������       �                     @        ^       a                   �p@�q�q�?             @       _       `                   0m@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        c       j                   @a@(N:!���?            �A@       d       i                 pff�?`2U0*��?             9@        e       f                    m@      �?              @       ������������������������       �                     @        g       h                   �_@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     1@        k       n                    `@�z�G��?             $@        l       m                     L@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        q       �                   �r@��R�(��?r            �e@       r       �                   �`@pIC'�T�?e            �b@       s       �                   P`@��(\���?7             T@       t       �                   8r@lGts��?%            �K@       u       ~                   `_@�:�]��?#            �I@       v       w                    �?���N8�?             E@       ������������������������       �                     B@        x       }                    �L@�q�q�?             @       y       z                    @K@�q�q�?             @        ������������������������       �                     �?        {       |                    `@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @               �                    �K@�<ݚ�?             "@       ������������������������       �                     @        �       �                    �L@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                     P@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     9@        �       �                    @K@:%�[��?.            �Q@       �       �                   @a@��S���?            �F@       �       �                   0d@X�<ݚ�?             B@        ������������������������       �                     @        �       �                    @C@��S���?             >@        �       �                   �]@�����H�?             "@        �       �                   �\@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �`@����X�?             5@       �       �                   @e@���y4F�?             3@        �       �                 033@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �a@      �?             0@        �       �                    @E@�<ݚ�?             "@        ������������������������       �                     �?        �       �                   �\@      �?              @        ������������������������       �                     @        �       �                   Pa@      �?             @        ������������������������       �                      @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                    �G@�����H�?             "@        ������������������������       �                     @        �       �                   �b@z�G�z�?             @        ������������������������       �                     @        �       �                    �I@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �a@8�Z$���?             :@        ������������������������       �                     $@        �       �                   b@      �?
             0@        ������������������������       �                      @        �       �                   �l@؇���X�?	             ,@        ������������������������       �                     @        �       �                    @L@      �?              @        ������������������������       �                     �?        �       �                   m@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    @I@�eP*L��?             6@        �       �                   �a@      �?              @        �       �                     G@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    @L@X�Cc�?             ,@        ������������������������       �                     @        �       �                     Q@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                    �E@�gtq���?S            �`@        �       �                   pb@ףp=
�?             $@        �       �                    @E@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                   0b@�<��S��?K            @_@        �       �                     H@ �q�q�?             8@        �       �                 `ff�?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     6@        �       �                    �?@VK��\�?>            @Y@        �       �                    i@� �	��?             9@        ������������������������       �                     @        �       �                    �O@�G�z��?             4@       �       �                 ����?ףp=
�?             $@       ������������������������       �                     @        �       �                    d@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     $@        �       �                    k@���=A�?0             S@        �       �                 ����?��.k���?             A@       �       �                    @N@��H�}�?             9@       �       �                    �?r�q��?             2@       �       �                    �?"pc�
�?             &@       ������������������������       �                      @        �       �                   �d@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                   �c@؇���X�?             @        ������������������������       �                     @        �       �                    �?      �?             @        ������������������������       �                      @        �       �                   @e@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �e@؇���X�?             @       ������������������������       �                     @        �       �                   Pa@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        �       �                   �c@d}h���?             E@       �       �                    �?�?�'�@�?             C@        �       �                    �?���Q��?             @       �       �                   `c@      �?             @        ������������������������       �                     �?        �       �                   �q@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �l@�C��2(�?            �@@        �       �                    @N@      �?              @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     9@        ������������������������       �                     @        �       �                    _@���c�H�?d            `b@        �       �                 033@XB���?+             M@       ������������������������       �        *             L@        ������������������������       �                      @        �                       ����?����?9            @V@                                 Xp@V������?            �B@                                b@8�Z$���?             :@                               �k@�X�<ݺ?             2@                                 ^@      �?              @                                �X@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     $@        	                          Q@      �?              @       
                         �L@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @                                 @L@���|���?             &@                               0`@      �?              @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @                                 y@4��?�?#             J@                             ����?HP�s��?!             I@                                �n@z�G�z�?             $@       ������������������������       �                      @        ������������������������       �                      @                                d@P���Q�?             D@       ������������������������       �                     A@                                 o@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @                                ��@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �t�bh�h)h,K ��h.��R�(KMKK��h^�B�  �5�;���?%e��?u��>P��?f�_O�?X驅���?O-�����?9��8���?�q�q�?_�_��?uPuP�?^Cy�5�?(������?�q�q�?�q�q�?�?�������?F]t�E�?]t�E�?              �?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?      �?              �?vb'vb'�?;�;��?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?        �u�y���?�).�u�?۳=۳=�?�0	�0	�?�������?���?      �?      �?��,d!�?��Moz��?              �?�������?�������?              �?�5��P�?(�����?      �?              �?      �?              �?      �?                      �?P?���O�?X`��?ffffff�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?        ����Ǐ�?����?      �?        ��<��<�?�a�a�?��y��y�?�a�a�?      �?        �q�q�?�q�q�?UUUUUU�?UUUUUU�?      �?              �?      �?      �?                      �?      �?              �?        'vb'vb�?�;�;�?a�|���?}���g�?              �?ȏ?~��?����?�;�;�?�؉�؉�?ffffff�?333333�?�������?333333�?              �?      �?              �?                      �?�������?UUUUUU�?X���oX�?��)A��?      �?        ��o��o�?�A�A�?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?�{����?�B!��?      �?        �m۶m��?�$I�$I�?      �?              �?      �?      �?                      �?333333�?�������?              �?      �?                      �?^N��)x�?����X�?�;����?W�+���?UUUUUU�?UUUUUU�?      �?        UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?              �?      �?                      �?|�W|�W�?�A�A�?���Q��?{�G�z�?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?        ffffff�?333333�?      �?      �?      �?                      �?      �?                      �?,�avp�?�*���}�?�Hs�9��?�-�q��?333333�?�������?�־a�?�<%�S��?�?}}}}}}�?�a�a�?��y��y�?              �?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?                      �?�q�q�?9��8���?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?      �?                      �?              �?�'�K=�?+l$Za�?�?�������?�q�q�?r�q��?              �?�?�������?�q�q�?�q�q�?      �?      �?              �?      �?                      �?�m۶m��?�$I�$I�?6��P^C�?(������?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?9��8���?�q�q�?              �?      �?      �?      �?              �?      �?      �?              �?      �?      �?                      �?      �?                      �?�q�q�?�q�q�?      �?        �������?�������?      �?              �?      �?              �?      �?        ;�;��?;�;��?              �?      �?      �?      �?        �$I�$I�?۶m۶m�?              �?      �?      �?      �?        �$I�$I�?۶m۶m�?      �?                      �?t�E]t�?]t�E�?      �?      �?      �?      �?              �?      �?              �?        �m۶m��?%I�$I��?              �?�m۶m��?�$I�$I�?      �?                      �?�\y@���?�Q�ߦ�?�������?�������?      �?      �?              �?      �?              �?        �l�����?�I+��?UUUUUU�?�������?      �?      �?              �?      �?                      �?:5r���?ce�F��?)\���(�?�Q����?              �?�������?�������?�������?�������?              �?      �?      �?              �?      �?              �?        �P^Cy�?��P^Cy�?�?�������?{�G�z�?
ףp=
�?�������?UUUUUU�?/�袋.�?F]t�E�?      �?        UUUUUU�?UUUUUU�?              �?      �?        ۶m۶m�?�$I�$I�?      �?              �?      �?      �?              �?      �?              �?      �?        �$I�$I�?۶m۶m�?              �?      �?      �?      �?                      �?              �?۶m۶m�?I�$I�$�?y�5���?������?�������?333333�?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?F]t�E�?]t�E�?      �?      �?              �?      �?                      �?      �?        /�����?4և����?�{a���?GX�i���?              �?      �?        e%+Y�J�?NmjS���?�g�`�|�?o0E>��?;�;��?;�;��?��8��8�?�q�q�?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?              �?              �?      �?�������?333333�?      �?                      �?      �?        F]t�E�?]t�E]�?      �?      �?              �?      �?                      �?ى�؉��?�N��N��?{�G�z�?q=
ףp�?�������?�������?              �?      �?        �������?ffffff�?              �?UUUUUU�?UUUUUU�?      �?                      �?      �?      �?      �?                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJF<KdhG        hNhG        hNhBKhDKhEh)h,K ��h.��R�(KK��h^�C              �?�t�bhQhchLC       ���R�hgKhhhkKh)h,K ��h.��R�(KK��hL�C       �t�bK��R�}�(hKhuMhvh)h,K ��h.��R�(KM��h}�B�D         �                    �?�#i����?�           ��@              �                   �a@�a�n��?l           ��@              h                    �?f	�B���?           0|@                                 @[@4և����?�            �q@                                   W@     ��?             @@        ������������������������       �                     $@                                   �G@8�A�0��?             6@        ������������������������       �                     @        	                          �`@�E��ӭ�?
             2@       
                           �N@������?	             1@                                 �X@؇���X�?             ,@        ������������������������       �                     @                                   Z@      �?              @                                  �K@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @                                ����?�q�q�?             @                                 �m@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?               g                   pe@��|,��?�             o@              :                    �G@Vβ���?�            @i@               9                    @G@����O��?+            �Q@              4                   Xq@.��<�?*            �P@              +                   �a@�2����?#            �K@               &                   `a@�X����?             6@              %                    �?@�0�!��?	             1@              $                    �?      �?             0@               !                   @_@8�Z$���?             *@        ������������������������       �                     @        "       #                    @F@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        '       *                    �?z�G�z�?             @       (       )                   o@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ,       3                   `i@�FVQ&�?            �@@        -       .                   �b@����X�?             @        ������������������������       �                     �?        /       2                    g@r�q��?             @        0       1                   pc@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     :@        5       6                   (r@�q�q�?             (@       ������������������������       �                     @        7       8                    @B@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ;       f                   Pe@tK���:�?V            ``@       <       e                    �R@8�Z$���?U            @`@       =       L                    @L@R��q�?T             `@       >       ?                    �H@@݈g>h�?2             S@        ������������������������       �        
             .@        @       A                   �j@Xny��?(            �N@        ������������������������       �                     :@        B       K                 ����?z�G�z�?            �A@       C       F                   k@6YE�t�?            �@@        D       E                   �`@���Q��?             @        ������������������������       �                     @        ������������������������       �                      @        G       H                   �q@@4և���?             <@       ������������������������       �                     5@        I       J                   �`@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        M       N                    [@�T`�[k�?"            �J@        ������������������������       �                     &@        O       T                   �\@����X�?             E@        P       S                    �M@      �?             @       Q       R                   l@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        U       d                    `P@�I�w�"�?             C@       V       ]                   P`@�z�G��?             >@        W       \                   �q@      �?
             $@       X       Y                 pff�?      �?              @        ������������������������       �                     @        Z       [                   `b@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        ^       _                   @c@z�G�z�?             4@       ������������������������       �                     $@        `       c                    �N@���Q��?             $@       a       b                   @f@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     G@        i       x                    �G@��U/��?q            `e@        j       w                    @��
P��?            �A@       k       l                   �[@�f7�z�?             =@        ������������������������       �                     @        m       n                    �?��+7��?             7@        ������������������������       �                     @        o       p                   �`@�q�q�?             2@        ������������������������       �                     @        q       r                    �@@؇���X�?             ,@        ������������������������       �                     �?        s       v                   �]@$�q-�?
             *@        t       u                   d@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     $@        ������������������������       �                     @        y       �                 `ff @      �?X             a@       z       �                    �Q@�w��#��?C             Y@       {       �                    �?     ��?A             X@       |       �                   �_@�99lMt�?2            �S@        }       �                    �P@      �?             @@       ~       �                   �k@П[;U��?             =@              �                   �^@D�n�3�?
             3@        ������������������������       �                     @        �       �                    �H@     ��?             0@        ������������������������       �                      @        �       �                   @b@d}h���?             ,@       ������������������������       �                     @        �       �                    �?և���X�?             @        ������������������������       �                      @        �       �                    @J@���Q��?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                    �?z�G�z�?             $@        �       �                 pff�?      �?             @        �       �                   �Z@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �\@r�q��?             @        ������������������������       �                      @        �       �                     J@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                 033�?��+7��?             G@       �       �                   (s@�<ݚ�?             B@       �       �                    �L@      �?             @@       �       �                    �?���y4F�?             3@        �       �                   �b@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   �_@d}h���?
             ,@        ������������������������       �                     @        �       �                   �d@      �?              @       �       �                   �`@      �?             @        �       �                    �J@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �k@      �?             @        ������������������������       �                     �?        �       �                    @K@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     *@        ������������������������       �                     @        �       �                    c@���Q��?             $@       �       �                    �?؇���X�?             @        ������������������������       �                     �?        �       �                    @J@r�q��?             @        ������������������������       �                     @        �       �                   �a@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �q@�����H�?             2@       ������������������������       �                     ,@        �       �                    @L@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     B@        �       �                   �w@
���n<�?M            �\@       �       �                    �?�Jl$G��?J            �[@       �       �                 `ff�?���y�?=            @V@        �       �                    �O@      �?             D@       �       �                    �?|��?���?             ;@        ������������������������       �                     @        �       �                   �l@�q�q�?             5@       �       �                   �\@      �?
             ,@        �       �                    @N@r�q��?             @        �       �                    @I@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �b@      �?              @       ������������������������       �                     @        �       �                    @L@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                   `p@8�Z$���?             *@        �       �                    �?���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        �       �                   �m@؇���X�?"            �H@       �       �                   0l@      �?             <@       �       �                    �?�C��2(�?             6@        ������������������������       �                     @        �       �                   �d@      �?
             0@       ������������������������       �        	             ,@        ������������������������       �                      @        �       �                   �a@r�q��?             @       ������������������������       �                     @        �       �                   �c@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     5@        �       �                    �?�eP*L��?             6@        �       �                   k@      �?              @       ������������������������       �                     @        �       �                   �]@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    S@X�Cc�?             ,@        �       �                   �b@և���X�?             @        ������������������������       �                     @        ������������������������       �                     @        �       �                   Pt@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    _@��s����?d             e@        ������������������������       �        )            �P@        �       �                   �f@�\�u��?;            �Y@        �       �                 ����?      �?              @       ������������������������       �                     @        ������������������������       �                     �?        �                         �b@V��N��?5            �W@       �                         �`@��UV�?)            �Q@       �       �                    @G@0G���ջ?              J@        ������������������������       �                     �?        �       �                    ^@`'�J�?            �I@        �       �                   Hp@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                     Q@`Ql�R�?            �G@       ������������������������       �                     E@        �                          `^@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?                              hff�?�����?	             3@        ������������������������       �                     @                                 n@@4և���?             ,@        ������������������������       �                      @                                c@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        	      
                   �?8����?             7@        ������������������������       �                     @                                 �G@b�2�tk�?	             2@        ������������������������       �                      @                                @n@     ��?             0@                               `\@      �?             $@        ������������������������       �                      @                                 �?      �?              @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �t�b��     h�h)h,K ��h.��R�(KMKK��h^�B0  �5�;���?%e��?���Ȇ�?ƿD\n��?�R�-���?AZ��@�?%I�$I��?n۶m۶�?      �?      �?              �?/�袋.�?颋.���?      �?        r�q��?�q�q�?�?xxxxxx�?�$I�$I�?۶m۶m�?              �?      �?      �?      �?      �?              �?      �?                      �?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?              �?        �RJ)���?���Zk��?z��~�X�?�&��? �
���?�]�����?IT�n��?o�Wc"=�?��7�}��?� O	��?�E]t��?]t�E]�?ZZZZZZ�?�������?      �?      �?;�;��?;�;��?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?�������?�������?      �?      �?      �?                      �?              �?>����?|���?�m۶m��?�$I�$I�?              �?�������?UUUUUU�?      �?      �?      �?                      �?      �?              �?        UUUUUU�?UUUUUU�?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?�T���?�����?;�;��?;�;��?Җ�%mI�?��-iK��?�P^Cy�?Cy�5��?      �?        C��6�S�?�}�K�`�?      �?        �������?�������?'�l��&�?e�M6�d�?�������?333333�?              �?      �?        n۶m۶�?�$I�$I�?      �?        �m۶m��?�$I�$I�?      �?                      �?              �?���!5��?"5�x+��?      �?        �m۶m��?�$I�$I�?      �?      �?UUUUUU�?UUUUUU�?              �?      �?                      �?����k�?�5��P�?ffffff�?333333�?      �?      �?      �?      �?              �?333333�?�������?      �?                      �?      �?        �������?�������?      �?        333333�?�������?۶m۶m�?�$I�$I�?              �?      �?                      �?      �?                      �?              �?      �?        g1��t�?Lg1��t�?_�_��?PuPu�?O#,�4��?a���{�?              �?zӛ����?Y�B��?      �?        UUUUUU�?UUUUUU�?              �?۶m۶m�?�$I�$I�?              �?�؉�؉�?;�;��?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?      �?      �?��(\���?��Q��?      �?      �?�o��o��?5H�4H��?      �?      �?��=���?�{a���?l(�����?(������?              �?      �?      �?              �?I�$I�$�?۶m۶m�?      �?        �$I�$I�?۶m۶m�?      �?        �������?333333�?      �?                      �?�������?�������?      �?      �?      �?      �?              �?      �?                      �?UUUUUU�?�������?              �?      �?      �?      �?                      �?      �?        Y�B��?zӛ����?�q�q�?9��8���?      �?      �?(������?6��P^C�?�������?�������?              �?      �?        ۶m۶m�?I�$I�$�?              �?      �?      �?      �?      �?      �?      �?              �?      �?              �?      �?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?      �?        �������?333333�?�$I�$I�?۶m۶m�?              �?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?              �?      �?              �?        �q�q�?�q�q�?              �?      �?      �?              �?      �?              �?                      �?�q�.�|�?<G�h���?镱��^�?5'��P�?p�\��?H?�я~�?      �?      �?{	�%���?	�%����?              �?UUUUUU�?UUUUUU�?      �?      �?UUUUUU�?�������?      �?      �?              �?      �?                      �?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?        ;�;��?;�;��?333333�?�������?      �?                      �?      �?        �$I�$I�?۶m۶m�?      �?      �?F]t�E�?]t�E�?              �?      �?      �?              �?      �?        �������?UUUUUU�?      �?              �?      �?              �?      �?                      �?t�E]t�?]t�E�?      �?      �?      �?              �?      �?              �?      �?        �m۶m��?%I�$I��?�$I�$I�?۶m۶m�?              �?      �?        �$I�$I�?۶m۶m�?              �?      �?                      �?�a�a�?z��y���?              �?�?�������?      �?      �?      �?                      �?��
br�?����F}�?6��9�?2~�ԓ��?�؉�؉�?vb'vb'�?      �?        �?�������?      �?      �?      �?                      �?W�+�ɕ?}g���Q�?              �?�������?�������?              �?      �?        ^Cy�5�?Q^Cy��?      �?        �$I�$I�?n۶m۶�?              �?UUUUUU�?�������?      �?                      �?d!Y�B�?8��Moz�?      �?        �8��8��?9��8���?              �?      �?      �?      �?      �?      �?              �?      �?              �?      �?              �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJؽ�hG        hNhG        hNhBKhDKhEh)h,K ��h.��R�(KK��h^�C              �?�t�bhQhchLC       ���R�hgKhhhkKh)h,K ��h.��R�(KK��hL�C       �t�bK��R�}�(hKhuMhvh)h,K ��h.��R�(KM��h}�B�G         �                 ����?�/�$�y�?�           ��@               �                    �?�mW��?�            �v@                                 @E@      �?�            �s@                                   п�z�G��?             >@        ������������������������       �                      @                                  ``@      �?             <@               
                    �F@      �?             0@               	                   �`@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     ,@                                hff�?      �?	             (@                                  �?      �?              @                                    Q@�q�q�?             @                               ����?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?                                   �P@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @               h                    @L@ظ�*���?�            �q@              O                   hq@���?�             l@              D                   �d@TL�n��?i            �f@              '                   �f@̌WZ�}�?I            �^@                                   �?      �?
             0@        ������������������������       �                      @               "                   �b@և���X�?	             ,@                                  �J@      �?              @       ������������������������       �                     @                !                   `_@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        #       $                 ������q�q�?             @        ������������������������       �                     �?        %       &                   `c@z�G�z�?             @        ������������������������       �                     @        ������������������������       �                     �?        (       =                   `@ܑ-Z���??            �Z@       )       8                   �o@H�ՠ&��?!             K@       *       7                    �?��S�ۿ?            �F@       +       6                   �d@�˹�m��?             C@       ,       5                   �a@@-�_ .�?            �B@        -       4                   k@      �?              @       .       /                   `Z@      �?             @        ������������������������       �                     �?        0       1                   �i@�q�q�?             @        ������������������������       �                     �?        2       3                   �_@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     =@        ������������������������       �                     �?        ������������������������       �                     @        9       :                    �C@X�<ݚ�?             "@        ������������������������       �                      @        ;       <                   d@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        >       ?                   Pk@�&=�w��?            �J@       ������������������������       �                     ;@        @       A                    _@$�q-�?             :@        ������������������������       �                     �?        B       C                 ����?`2U0*��?             9@       ������������������������       �                     8@        ������������������������       �                     �?        E       L                   �b@���#�İ?             �M@       F       G                   `a@0�)AU��?            �L@       ������������������������       �                    �G@        H       K                    b@ףp=
�?             $@       I       J                    �B@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        M       N                    �E@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        P       ]                   @c@��V#�?            �E@        Q       X                   �`@�\��N��?             3@       R       W                   (@"pc�
�?             &@       S       T                    �?ףp=
�?             $@       ������������������������       �                      @        U       V                   `c@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        Y       Z                   0a@      �?              @        ������������������������       �                     @        [       \                     J@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ^       g                 ����?�q�q�?             8@       _       f                   @r@�GN�z�?             6@        `       a                    �C@r�q��?             @        ������������������������       �                     @        b       c                    �?�q�q�?             @        ������������������������       �                     �?        d       e                   @_@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �        	             0@        ������������������������       �                      @        i       �                    �P@D�n�3�?'            �L@       j       w                   �k@�`���?$            �H@        k       v                 833�?������?             1@       l       u                     P@�q�q�?	             (@       m       t                    @N@���!pc�?             &@       n       o                   @Z@և���X�?             @        ������������������������       �                      @        p       s                   b@���Q��?             @       q       r                   �i@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        x       �                   �u@      �?             @@       y       z                   @`@�q�q�?             >@        ������������������������       �                     @        {       �                   p`@\X��t�?             7@        |       }                   �Z@���!pc�?             &@        ������������������������       �                     �?        ~       �                 @33�?z�G�z�?             $@               �                   �d@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                   pa@�q�q�?
             (@        ������������������������       �                     @        �       �                   �c@      �?              @       �       �                    �N@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                      @        �       �                    �?J��D��?&             K@        �       �                   �h@"pc�
�?             &@        ������������������������       �                     @        �       �                   �`@      �?             @       ������������������������       �                      @        ������������������������       �                      @        �       �                 833�?8�$�>�?             �E@       �       �                   `o@������?             A@       �       �                    迴C��2(�?             6@        ������������������������       �                     �?        �       �                     G@�����?             5@        �       �                    @E@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?      �?             0@       �       �                   @V@ףp=
�?             $@        ������������������������       �                     @        �       �                   �_@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                   8p@      �?	             (@        ������������������������       �                     @        �       �                    �?�q�q�?             "@       �       �                   �p@      �?             @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                 ����?�<ݚ�?             "@       �       �                   �O@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �L@     ��?�             w@       �       �                 033�?�q�qT�?{             h@        �       �                   (s@�U���?*             O@       �       �                   �b@�q�q�?%             K@       �       �                    �?z�G�z�?             D@       �       �                   �]@     ��?             @@        ������������������������       �                     &@        �       �                 ����?�q�q�?             5@       �       �                    �F@     ��?             0@        ������������������������       �                     @        �       �                   �m@���|���?             &@        �       �                   �`@���Q��?             @       �       �                    @K@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   �`@r�q��?             @        ������������������������       �                     @        �       �                   �a@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                   �g@d}h���?             ,@        ������������������������       �                      @        �       �                   �d@�8��8��?
             (@       ������������������������       �                     @        �       �                   �i@r�q��?             @        ������������������������       �                     @        �       �                    l@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                     J@      �?              @        ������������������������       �                     @        �       �                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   �g@�����D�?Q            @`@        ������������������������       �                     A@        �       �                   �c@      �?<             X@       �       �                   �a@�+ت�M�?1            �S@       �       �                   �Z@�����?"            �H@        ������������������������       �                     �?        �       �                    �J@     ��?!             H@        �       �                   �a@8����?             7@       �       �                    ]@@�0�!��?             1@        �       �                   m@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        	             *@        �       �                   �c@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                   @_@HP�s��?             9@       ������������������������       �        
             .@        �       �                    _@z�G�z�?             $@        �       �                 033@���Q��?             @       �       �                   @a@�q�q�?             @        ������������������������       �                     �?        �       �                   �o@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     >@        �       �                    @@�0�!��?             1@       �       �                   �e@�r����?	             .@       ������������������������       �                     *@        ������������������������       �                      @        �       �                   �e@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �                         �z@�Ra����?o             f@       �                       ���@ܷ��?��?m            �e@       �                          �?x�c/y[�?T            �`@       �       �                   @\@��r._�?3            �T@        ������������������������       �                     =@        �       	                   c@Ȩ�I��?"            �J@       �                         P`@fP*L��?             F@        �       �                   �\@      �?	             (@        ������������������������       �                     @        �       �                    @O@؇���X�?             @       ������������������������       �                     @                                  `P@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?                                 �?      �?             @@                               pb@�IєX�?             1@       ������������������������       �        	             *@                              `ff�?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     .@        
                        `a@�<ݚ�?             "@       ������������������������       �                     @                                 �?      �?             @        ������������������������       �                      @        ������������������������       �                      @                                �[@0G���ջ?!             J@        ������������������������       �        
             2@                                 �R@l��\��?             A@                             ����?      �?             @@                                `c@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     ;@        ������������������������       �                      @                                  P@�(\����?             D@       ������������������������       �                     ?@                                �]@�����H�?             "@                                �[@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �t�bh�h)h,K ��h.��R�(KMKK��h^�B�  L�f���?Z�L��?J�=���?l�g��?      �?      �?333333�?ffffff�?      �?              �?      �?      �?      �?      �?      �?      �?                      �?              �?      �?      �?      �?      �?UUUUUU�?UUUUUU�?      �?      �?              �?      �?              �?        �������?�������?      �?                      �?              �?&W�+��?g���Q��?O贁N�?ƒ_,���?�ʨ�ʨ�?�������?�[<�œ�?����?      �?      �?              �?�$I�$I�?۶m۶m�?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?UUUUUU�?      �?        �������?�������?              �?      �?        ��	�N�?�rp�_��?������?{	�%���?�������?�?��P^Cy�?^Cy�5�?S�n0E�?к����?      �?      �?      �?      �?              �?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?              �?              �?                      �?      �?        r�q��?�q�q�?              �?�m۶m��?�$I�$I�?      �?                      �?tHM0���?�x+�R�?      �?        �؉�؉�?;�;��?              �?���Q��?{�G�z�?      �?                      �?��N��?'u_[�?��Gp�?p�}��?      �?        �������?�������?�������?UUUUUU�?              �?      �?              �?              �?      �?              �?      �?        eMYS֔�?6eMYS��?y�5���?�5��P�?/�袋.�?F]t�E�?�������?�������?      �?              �?      �?              �?      �?                      �?      �?      �?              �?      �?      �?              �?      �?        UUUUUU�?�������?�袋.��?]t�E�?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?              �?              �?        l(�����?(������?����S�?և���X�?xxxxxx�?�?UUUUUU�?UUUUUU�?F]t�E�?t�E]t�?�$I�$I�?۶m۶m�?      �?        �������?333333�?      �?      �?              �?      �?              �?              �?                      �?      �?              �?      �?UUUUUU�?UUUUUU�?              �?��Moz��?!Y�B�?t�E]t�?F]t�E�?      �?        �������?�������?      �?      �?      �?                      �?              �?�������?�������?      �?              �?      �?      �?      �?              �?      �?                      �?      �?              �?        _B{	�%�?�^B{	��?F]t�E�?/�袋.�?              �?      �?      �?              �?      �?        �5eMYS�?6eMYS��?�?xxxxxx�?F]t�E�?]t�E�?              �?�a�a�?=��<���?�������?�������?              �?      �?              �?      �?�������?�������?              �?�������?�������?      �?                      �?              �?      �?      �?      �?        UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?9��8���?�q�q�?      �?      �?              �?      �?                      �?      �?      �?UUUUUU�?UUUUU��?�9�s��?c�1��?UUUUUU�?UUUUUU�?ffffff�?ffffff�?      �?      �?              �?UUUUUU�?UUUUUU�?      �?      �?              �?]t�E]�?F]t�E�?�������?333333�?UUUUUU�?UUUUUU�?      �?                      �?              �?�������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?              �?I�$I�$�?۶m۶m�?              �?UUUUUU�?UUUUUU�?      �?        �������?UUUUUU�?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?      �?      �?        �������?�������?      �?                      �?z�z��?z�z��?              �?      �?      �?h *�3�?�w��	��?����X�?^N��)x�?      �?              �?      �?8��Moz�?d!Y�B�?�������?ZZZZZZ�?      �?      �?              �?      �?                      �?UUUUUU�?UUUUUU�?      �?                      �?{�G�z�?q=
ףp�?              �?�������?�������?�������?333333�?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?                      �?              �?              �?ZZZZZZ�?�������?�������?�?      �?                      �?      �?      �?              �?      �?        ]t�E�?]t�E]�?a���{�?��=���?o�Wc"=�?�*g���?ە�]���?�ڕ�]��?              �?�	�[���?+�R��?]t�E]�?颋.���?      �?      �?              �?۶m۶m�?�$I�$I�?      �?              �?      �?              �?      �?              �?      �?�?�?              �?      �?      �?      �?                      �?              �?9��8���?�q�q�?      �?              �?      �?              �?      �?        �؉�؉�?vb'vb'�?              �?�������?------�?      �?      �?�������?�������?      �?                      �?              �?      �?        �������?333333�?              �?�q�q�?�q�q�?      �?      �?              �?      �?                      �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJX��vhG        hNhG        hNhBKhDKhEh)h,K ��h.��R�(KK��h^�C              �?�t�bhQhchLC       ���R�hgKhhhkKh)h,K ��h.��R�(KK��hL�C       �t�bK��R�}�(hKhuMhvh)h,K ��h.��R�(KM��h}�B@D         �                 ����?���
%�?�           ��@               �                    �?���u�J�?�            �v@              b                    @M@�{�Mk��?�            Ps@                                 �P@>�b@��?�            �o@               
                    �?؇���X�?             ,@              	                   �[@"pc�
�?	             &@                                 �Z@�q�q�?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @               G                   q@��[�-�?�            �m@                                   �F@��zi��?o            �f@                                  �d@xL��N�?1            �R@        ������������������������       �                     =@                                   �B@��S�ۿ?            �F@        ������������������������       �        	             &@                                   �?l��\��?             A@                                 �d@��a�n`�?             ?@        ������������������������       �                     �?                                  l@��S�ۿ?             >@                                   �?؇���X�?	             ,@                                   j@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                   @D@�C��2(�?             &@                                  `j@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        	             0@        ������������������������       �                     @        !       2                   �_@r�i�+$�?>             [@        "       -                    @K@��.k���?             A@       #       ,                    �?���N8�?
             5@       $       %                   @Z@�S����?             3@        ������������������������       �                     �?        &       +                    �J@�����H�?             2@       '       (                    �?r�q��?             (@        ������������������������       �                     �?        )       *                   �a@�C��2(�?             &@       ������������������������       �                     $@        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        .       /                   @Z@8�Z$���?             *@        ������������������������       �                     @        0       1                   �i@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        3       :                   �l@�x
�2�?-            �R@       4       5                    �L@�(\����?             D@       ������������������������       �                    �B@        6       9                 @33�?�q�q�?             @       7       8                   �h@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ;       <                   �l@�t����?             A@        ������������������������       �                      @        =       D                    @J@      �?             @@       >       C                   �p@     ��?             0@       ?       @                    �?�q�q�?	             (@        ������������������������       �                     @        A       B                   �l@�<ݚ�?             "@        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        E       F                   �a@      �?	             0@        ������������������������       �                     �?        ������������������������       �                     .@        H       a                    �L@�����?"            �L@       I       V                    �H@�1�`jg�?!            �K@       J       O                   8r@*;L]n�?             >@        K       N                   hq@8�Z$���?             *@        L       M                   �_@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     "@        P       Q                   �a@�t����?             1@       ������������������������       �                     &@        R       U                   �c@�q�q�?             @        S       T                   Pa@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        W       \                    �?H%u��?             9@        X       Y                   ``@      �?              @        ������������������������       �                     �?        Z       [                   r@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ]       `                    @K@�IєX�?
             1@       ^       _                   �r@�C��2(�?             &@        ������������������������       �                     �?        ������������������������       �                     $@        ������������������������       �                     @        ������������������������       �                      @        c       �                   Pd@���>4��?&             L@       d       }                     Q@j���� �?"            �I@       e       |                   �a@�X���?             F@       f       g                    �?�Gi����?            �B@        ������������������������       �                      @        h       s                   P`@l��[B��?             =@        i       r                   �`@�q�q�?             .@       j       o                    �?�θ�?             *@       k       n                 hff�?�����H�?             "@       l       m                 ����?      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        p       q                   @_@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                      @        t       {                 ����?����X�?
             ,@       u       v                    �N@X�<ݚ�?             "@        ������������������������       �                     @        w       z                   �]@z�G�z�?             @        x       y                    X@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ~                          c@؇���X�?             @       ������������������������       �                     @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �O@�	j*D�?%             J@        ������������������������       �                     6@        �       �                    �L@��S���?             >@       �       �                   �Z@z�G�z�?             .@        ������������������������       �                     �?        �       �                   n@؇���X�?             ,@        ������������������������       �                     @        �       �                   �d@����X�?             @        ������������������������       �                     @        �       �                    �G@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                   0j@������?	             .@        �       �                 hff�?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        �       �                    �?r�q��?             (@       �       �                    p@���Q��?             @       �       �                    �Q@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        �       �                 pff�?|��T+[�?�            Pw@        �       �                   �_@<�\`*��?9             U@       �       �                    �H@��|�5��?!            �G@        ������������������������       �                     &@        �       �                   �`@<ݚ)�?             B@        �       �                   @\@�\��N��?             3@        ������������������������       �                     @        �       �                     O@����X�?
             ,@       �       �                 `ff�?�θ�?	             *@        ������������������������       �                     �?        �       �                    @L@r�q��?             (@        �       �                    �I@�q�q�?             @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �       �                   �a@�IєX�?             1@        �       �                    �Q@      �?              @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     "@        �       �                    �?��+��?            �B@        ������������������������       �                     @        �       �                   0a@��.k���?             A@        ������������������������       �                     @        �       �                   �f@��S���?             >@        ������������������������       �                     @        �       �                   Pi@�û��|�?             7@        �       �                   �\@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        �       �                   �j@      �?             0@        ������������������������       �                     @        �       �                   0c@���!pc�?	             &@       �       �                   �a@      �?             @       �       �                    �?���Q��?             @       �       �                   @`@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                 `ff @^�R|���?�            r@       �       �                   P`@@�G��S�?}            @i@        �       �                   �c@�VM�?3            @V@       �       �                    �P@�I�w�"�?+             S@       �       �                   �]@���@��?)            �R@        ������������������������       �                     6@        �       �                   �m@�	j*D�?             J@       �       �                   p`@     ��?             @@       �       �                    @O@�GN�z�?
             6@       �       �                 033�?�KM�]�?	             3@        �       �                 ����?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     0@        ������������������������       �                     @        �       �                    �?z�G�z�?             $@       �       �                    �F@���Q��?             @        ������������������������       �                     �?        �       �                   �V@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        �       �                   �b@R���Q�?
             4@       ������������������������       �                     (@        �       �                   �p@      �?              @       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        �       �                   `l@8�Z$���?             *@       ������������������������       �                      @        �       �                   �z@���Q��?             @       ������������������������       �                      @        ������������������������       �                     @        �       �                   0s@h��)�~�?J            @\@       �       �                    �M@b �57�?C            �Y@       �       �                    c@H%u��?#             I@       �       �                   `k@�Ń��̧?             E@       �       �                   �j@���N8�?             5@       ������������������������       �                     3@        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     5@        �       �                   �e@      �?              @       �       �                 ����?����X�?             @        �       �                    �G@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     �?        �       �                     Q@�O4R���?             �J@       ������������������������       �                     A@        �       �                   �b@�}�+r��?             3@       ������������������������       �        
             2@        ������������������������       �                     �?        �       �                   �s@���Q��?             $@        ������������������������       �                     @        ������������������������       �                     @        �                         �l@X��%�?4            �U@                                 �?,���i�?            �D@                               pb@�#-���?            �A@                               @b@ ��WV�?             :@       ������������������������       �                     5@                                �b@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @              
                   �?�<ݚ�?             "@             	                    P@      �?              @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     �?                                �`@�q�q�?             @                                @e@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     G@        �t�bh�h)h,K ��h.��R�(KMKK��h^�B  ��\���?��Q���?�r�z[��?=�
I��?o�:�x�?�![��?k�Dly(�?S��N^�?�$I�$I�?۶m۶m�?F]t�E�?/�袋.�?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?,��E1N�?P���:��?��_��_�?h�h��?>�S��?L�Ϻ��?      �?        �������?�?      �?        ------�?�������?�s�9��?�c�1Ƹ?              �?�������?�?۶m۶m�?�$I�$I�?UUUUUU�?UUUUUU�?              �?      �?        ]t�E�?F]t�E�?      �?      �?      �?                      �?      �?              �?              �?        ���Kh�?��Kh/�?�?�������?��y��y�?�a�a�?^Cy�5�?(������?      �?        �q�q�?�q�q�?UUUUUU�?�������?      �?        F]t�E�?]t�E�?              �?      �?                      �?      �?        ;�;��?;�;��?      �?        �m۶m��?�$I�$I�?              �?      �?        �n0E>�?o0E>��?333333�?�������?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?        �������?�������?              �?      �?      �?      �?      �?�������?�������?      �?        �q�q�?9��8���?      �?                      �?      �?              �?      �?              �?      �?        Q^Cy��?^Cy�5�?��k߰�?��)A��?""""""�?�������?;�;��?;�;��?      �?      �?              �?      �?                      �?<<<<<<�?�?      �?        UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?        )\���(�?���Q��?      �?      �?              �?۶m۶m�?�$I�$I�?              �?      �?        �?�?]t�E�?F]t�E�?              �?      �?              �?                      �?n۶m۶�?I�$I�$�?ZZZZZZ�?�������?�E]t��?]t�E�?#�u�)��?o0E>��?              �?���=��?GX�i���?UUUUUU�?UUUUUU�?�؉�؉�?ى�؉��?�q�q�?�q�q�?      �?      �?              �?      �?                      �?      �?      �?      �?                      �?      �?        �m۶m��?�$I�$I�?r�q��?�q�q�?      �?        �������?�������?      �?      �?              �?      �?                      �?      �?                      �?۶m۶m�?�$I�$I�?      �?              �?      �?              �?      �?              �?        ;�;��?vb'vb'�?              �?�?�������?�������?�������?              �?۶m۶m�?�$I�$I�?      �?        �m۶m��?�$I�$I�?      �?              �?      �?              �?      �?        �?wwwwww�?UUUUUU�?UUUUUU�?      �?                      �?UUUUUU�?�������?�������?333333�?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?+�O��d�?��Ǧ�?�a�a�?=��<���?x6�;��?br1���?              �?�8��8��?��8��8�?y�5���?�5��P�?              �?�m۶m��?�$I�$I�?ى�؉��?�؉�؉�?              �?�������?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?�?�?      �?      �?              �?      �?                      �?*�Y7�"�?�S�n�?              �?�������?�?      �?        �������?�?              �?8��Moz�?��,d!�?۶m۶m�?�$I�$I�?              �?      �?              �?      �?              �?F]t�E�?t�E]t�?      �?      �?333333�?�������?      �?      �?      �?                      �?              �?              �?      �?        �W��H��?�@�m�?z��~�X�?�Q`ҩ�?NmjS���?Y�JV���?�5��P�?����k�?к����?L�Ϻ��?              �?;�;��?vb'vb'�?      �?      �?]t�E�?�袋.��?(�����?�k(���?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?        �������?�������?333333�?�������?              �?      �?      �?              �?      �?              �?        333333�?333333�?              �?      �?      �?              �?      �?              �?        ;�;��?;�;��?      �?        333333�?�������?              �?      �?        Ź�Q��?�(�u���?�H%�e�?��VC��?���Q��?)\���(�?�a�a�?��<��<�?�a�a�?��y��y�?              �?      �?      �?              �?      �?                      �?      �?      �?�m۶m��?�$I�$I�?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?�x+�R�?:�&oe�?              �?(�����?�5��P�?              �?      �?        �������?333333�?      �?                      �?��֡�l�? ��2)�?8��18�?�����?_�_�?�A�A�?;�;��?O��N���?              �?�������?�������?      �?                      �?�q�q�?9��8���?      �?      �?              �?      �?                      �?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ���EhG        hNhG        hNhBKhDKhEh)h,K ��h.��R�(KK��h^�C              �?�t�bhQhchLC       ���R�hgKhhhkKh)h,K ��h.��R�(KK��hL�C       �t�bK��R�}�(hKhuM'hvh)h,K ��h.��R�(KM'��h}�B�I         D                    �G@�r,��?�           ��@               =                    �?��bu<	�?q            `f@              $                   �c@r�u���?h            �d@                                  `a@�p ��?2            �T@                                 @q@�G\�c�?'            @P@                                 �]@�2�o�U�?!            �K@                                   \@8�A�0��?             6@        ������������������������       �                     @        	       
                   �h@������?
             1@        ������������������������       �                     @                                ����?���Q��?             $@        ������������������������       �                      @                                   �?      �?              @        ������������������������       �                     �?                                   �F@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?                                   �?<���D�?            �@@                                  @j@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                  �`@ףp=
�?             >@                                   �?�z�G��?             $@       ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     4@        ������������������������       �                     $@               #                   `a@������?             1@              "                    @G@�q�q�?             (@              !                    �?���Q��?             $@                                  �Y@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @        %       ,                   �[@�m(�X�?6            @U@        &       )                    @C@և���X�?             @        '       (                   �e@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        *       +                    �?      �?             @        ������������������������       �                     �?        ������������������������       �                     @        -       <                    @D@�7��?0            �S@        .       5                   `e@(N:!���?            �A@        /       0                    �A@      �?             (@        ������������������������       �                     @        1       4                   �d@      �?             @       2       3                    @B@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        6       7                    �C@�nkK�?             7@       ������������������������       �                     0@        8       ;                   �l@؇���X�?             @        9       :                 `ff�?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                    �E@        >       C                    �?�8��8��?	             (@       ?       B                   �_@ףp=
�?             $@        @       A                   @a@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        E       d                   @E@v�1>'��?_           X�@        F       G                   �\@P>�7���?D            @]@        ������������������������       �                     E@        H       c                    �?b����o�?.            �R@       I       R                 033�?)O���?             B@        J       Q                   �c@      �?
             (@       K       L                    �?"pc�
�?	             &@        ������������������������       �                     �?        M       N                   �`@ףp=
�?             $@        ������������������������       �                     @        O       P                   a@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        S       \                    �?�q�q�?             8@       T       Y                   �a@؇���X�?
             ,@       U       V                   P`@�8��8��?             (@       ������������������������       �                     @        W       X                    �?z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        Z       [                   �b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ]       ^                   �]@���Q��?             $@        ������������������������       �                      @        _       `                     K@      �?              @        ������������������������       �                     �?        a       b                    �O@؇���X�?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                    �C@        e       �                   �`@T]�z�?           `{@        f       �                   ``@įDg50�?�            @i@        g       �                 033�?*-ڋ�p�?7            @S@       h       o                   @i@      �?(             M@        i       j                   �[@"pc�
�?	             &@        ������������������������       �                     @        k       l                   `^@����X�?             @        ������������������������       �                     �?        m       n                 @33�?r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @        p       u                    ]@�[�IJ�?            �G@        q       t                 ����?�8��8��?             (@        r       s                   @Z@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        v       �                 033�?�xGZ���?            �A@       w       �                   �]@���@M^�?             ?@       x       }                   �X@      �?             4@        y       |                    �?r�q��?             @       z       {                   �m@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        ~                           �I@X�Cc�?
             ,@        ������������������������       �                      @        �       �                    �?      �?             (@        ������������������������       �                      @        �       �                   @^@ףp=
�?             $@        �       �                   �l@z�G�z�?             @        ������������������������       �                     �?        �       �                    �J@      �?             @        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?"pc�
�?             &@        �       �                    @Q@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?�}�+r��?             3@       ������������������������       �                     1@        �       �                   �\@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    @K@L.��:��?P            @_@        �       �                    `@����X�?             <@       �       �                    �I@r�q��?             8@        �       �                    �?�θ�?             *@       �       �                   �p@r�q��?             (@       �       �                   �^@      �?              @       �       �                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     �?        �       �                    �?�C��2(�?             &@        �       �                   �f@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     "@        ������������������������       �                     @        �       �                 833�?�^'�ë�?=            @X@        �       �                    �?      �?             ,@       �       �                    @O@�q�q�?	             (@       �       �                   `n@      �?              @        ������������������������       �                     @        �       �                    �?�q�q�?             @        ������������������������       �                     �?        �       �                   �q@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    �P@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �       �                   0l@P��BNֱ?2            �T@        ������������������������       �                     A@        �       �                 `ff@��<D�m�?            �H@       �       �                   `_@�?�|�?            �B@       ������������������������       �                     =@        �       �                   �_@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    n@r�q��?             (@        ������������������������       �                      @        ������������������������       �                     $@        �       �                    �L@�Zc!J��?�            �m@       �       �                 ����?���qK�?Y            �`@       �       �                   �q@,sI�v�?;            �V@       �       �                 ����?���Lͩ�?1            �R@       �       �                    �?�F��O�?/            @R@       �       �                   `@ �Cc}�?$             L@       �       �                   �l@�>4և��?             <@        �       �                   �\@�n_Y�K�?
             *@        ������������������������       �                     @        �       �                   �j@X�<ݚ�?             "@       �       �                   �^@�q�q�?             @       �       �                   �`@���Q��?             @        ������������������������       �                      @        �       �                   �h@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �        
             .@        �       �                    @I@h�����?             <@        �       �                   �p@      �?              @       �       �                   �m@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     4@        ������������������������       �                     1@        �       �                    �J@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �f@������?
             .@       �       �                   `c@d}h���?	             ,@        �       �                   �r@      �?             @        ������������������������       �                      @        �       �                   t@      �?             @        ������������������������       �                      @        �       �                    �?      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        �       �                   �h@�^�����?            �E@        �       �                     J@���|���?             &@        ������������������������       �                     @        ������������������������       �                     @        �       �                    �?     ��?             @@        �       �                   �u@���Q��?             @       ������������������������       �                      @        ������������������������       �                     @        �       �                   c@PN��T'�?             ;@       �       �                   @b@"pc�
�?             6@       �       �                 ����?؇���X�?             5@        ������������������������       �                     $@        �       �                    �?���!pc�?	             &@       �       �                   �a@      �?              @        ������������������������       �                     @        �       �                    @���Q��?             @       �       �                   �d@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        �                       ����?\x�R:��?;            �Y@                                �c@���!pc�?$            �P@                               �_@؇���X�?            �A@        ������������������������       �                     1@                                 �?�E��ӭ�?             2@                             ����?     ��?             0@                               �g@���!pc�?             &@        ������������������������       �                     @              
                   �N@և���X�?             @              	                  Pb@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                      @                                pe@�P�*�?             ?@                                n@r�q��?             8@                             ����?�	j*D�?             *@                               Pd@"pc�
�?             &@                               0a@�q�q�?             @        ������������������������       �                     @                                 @M@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                      @                                �Z@"pc�
�?             &@        ������������������������       �                      @        ������������������������       �                     "@        ������������������������       �                     @                                �a@�L���?            �B@        ������������������������       �                     &@                                  b@ȵHPS!�?             :@        ������������������������       �                     �?        !      &                   �?HP�s��?             9@       "      %                033�?ףp=
�?             4@        #      $                  xu@���Q��?             @       ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     .@        ������������������������       �                     @        �t�b���      h�h)h,K ��h.��R�(KM'KK��h^�Bp  �292ȯ�?�f����?��e㛡�?��49ȼ�?E���w��?v���?dp>�c�?8��18�?S+�R+��?[��Z���?־a��?�S�<%��?/�袋.�?颋.���?      �?        �?xxxxxx�?              �?�������?333333�?      �?              �?      �?      �?        �$I�$I�?۶m۶m�?              �?      �?        |���?|���?UUUUUU�?UUUUUU�?              �?      �?        �������?�������?ffffff�?333333�?      �?                      �?      �?                      �?�?xxxxxx�?UUUUUU�?UUUUUU�?�������?333333�?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?              �?]]]]]]�?�?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?              �?      �?              �?      �?              �?      �?        ��[��[�?�A�A�?|�W|�W�?�A�A�?      �?      �?      �?              �?      �?      �?      �?              �?      �?                      �?�Mozӛ�?d!Y�B�?      �?        ۶m۶m�?�$I�$I�?      �?      �?              �?      �?              �?              �?        UUUUUU�?UUUUUU�?�������?�������?      �?      �?              �?      �?                      �?              �?�AVO��?@�T��?�)��)��?��Y��Y�?              �?�6�i�?�X�%��?��8��8�?9��8���?      �?      �?/�袋.�?F]t�E�?              �?�������?�������?      �?        �������?�������?              �?      �?                      �?UUUUUU�?UUUUUU�?�$I�$I�?۶m۶m�?UUUUUU�?UUUUUU�?              �?�������?�������?              �?      �?              �?      �?      �?                      �?333333�?�������?              �?      �?      �?              �?۶m۶m�?�$I�$I�?      �?                      �?              �?��'����?� 산�?�F�tj�?B���be�?��cj`��??!��O��?      �?      �?/�袋.�?F]t�E�?      �?        �m۶m��?�$I�$I�?              �?�������?UUUUUU�?              �?      �?        m�w6�;�?���
b�?UUUUUU�?UUUUUU�?      �?      �?      �?                      �?              �?�_�_�?�A�A�?�s�9��?�c�1��?      �?      �?�������?UUUUUU�?      �?      �?      �?                      �?      �?        �m۶m��?%I�$I��?      �?              �?      �?      �?        �������?�������?�������?�������?              �?      �?      �?              �?      �?                      �?/�袋.�?F]t�E�?      �?      �?              �?      �?              �?                      �?(�����?�5��P�?              �?      �?      �?      �?                      �?;�O��n�?1�Zd�?�$I�$I�?�m۶m��?UUUUUU�?�������?�؉�؉�?ى�؉��?UUUUUU�?�������?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?              �?              �?      �?        F]t�E�?]t�E�?      �?      �?              �?      �?                      �?      �?        ���Id�?=�L�v��?      �?      �?�������?�������?      �?      �?      �?        UUUUUU�?UUUUUU�?              �?      �?      �?              �?      �?              �?      �?              �?      �?                      �?���ˊ��?��FS���?              �?և���X�?��S�r
�?к����?*�Y7�"�?              �?      �?      �?      �?                      �?UUUUUU�?�������?      �?                      �?����c�?�<�"h8�?*b���"�?�;��?l�l��?��I��I�?�6�i�?�K~��?�իW�^�?�P�B�
�?%I�$I��?۶m۶m�?�$I�$I�?�m۶m��?;�;��?ى�؉��?      �?        �q�q�?r�q��?UUUUUU�?UUUUUU�?333333�?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?                      �?      �?        �m۶m��?�$I�$I�?      �?      �?      �?      �?      �?                      �?      �?              �?              �?              �?      �?              �?      �?        wwwwww�?�?I�$I�$�?۶m۶m�?      �?      �?              �?      �?      �?      �?              �?      �?      �?                      �?      �?                      �?֔5eMY�?�5eMYS�?]t�E]�?F]t�E�?              �?      �?              �?      �?�������?333333�?      �?                      �?h/�����?&���^B�?F]t�E�?/�袋.�?�$I�$I�?۶m۶m�?              �?t�E]t�?F]t�E�?      �?      �?              �?333333�?�������?      �?      �?      �?                      �?              �?              �?      �?                      �?\mMw��?R�yY�'�?F]t�E�?t�E]t�?۶m۶m�?�$I�$I�?      �?        �q�q�?r�q��?      �?      �?F]t�E�?t�E]t�?      �?        �$I�$I�?۶m۶m�?      �?      �?              �?      �?              �?              �?                      �?�RJ)���?�Zk����?UUUUUU�?UUUUUU�?vb'vb'�?;�;��?/�袋.�?F]t�E�?UUUUUU�?UUUUUU�?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?F]t�E�?/�袋.�?      �?                      �?      �?        L�Ϻ��?}���g�?              �?�؉�؉�?��N��N�?      �?        {�G�z�?q=
ףp�?�������?�������?�������?333333�?              �?      �?                      �?              �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ:9)bhG        hNhG        hNhBKhDKhEh)h,K ��h.��R�(KK��h^�C              �?�t�bhQhchLC       ���R�hgKhhhkKh)h,K ��h.��R�(KK��hL�C       �t�bK��R�}�(hKhuMhvh)h,K ��h.��R�(KM��h}�B�D         �                    @K@T8���?�           ��@              _                 ����?����_�?�             x@                                  I@d�K��?�            @n@                                  @\@PN��T'�?             ;@               
                    �?�	j*D�?             *@                                 �Z@      �?             (@       ������������������������       �                      @               	                    @I@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     ,@               @                   �c@RB)��.�?�            �j@                                  �]@t�I��n�?A            @]@                                  @[@��
ц��?             :@        ������������������������       �                      @                                   @G@�q�q�?
             2@                                  @E@8�Z$���?             *@                                  �\@����X�?             @                                 �a@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @                                   �?z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @               ?                 ����?|�H���?1            �V@              "                    @E@z\�3�?,            �S@               !                    `@�nkK�?             7@                                   `_@�����H�?             "@       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     ,@        #       ,                   `a@������?              L@        $       +                   r@�q�q�?             8@       %       *                   �`@�㙢�c�?             7@       &       )                   �\@�	j*D�?             *@        '       (                   �l@      �?              @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     $@        ������������������������       �                     �?        -       8                   Hp@     ��?             @@       .       7                   �k@�KM�]�?             3@        /       6                    �?����X�?             @       0       1                    �I@���Q��?             @        ������������������������       �                      @        2       5                    b@�q�q�?             @       3       4                   �^@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     (@        9       >                    �G@$�q-�?             *@        :       ;                   �_@z�G�z�?             @        ������������������������       �                     @        <       =                   0b@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     (@        A       ^                    r@H;T*St�?A            �X@       B       ]                    �?z���=��?3            @S@       C       X                   Hq@F.< ?�?-            �P@       D       I                   �[@Riv����?)             M@        E       F                   @[@X�<ݚ�?             "@        ������������������������       �                      @        G       H                    @G@����X�?             @        ������������������������       �                     @        ������������������������       �                      @        J       K                   pk@Hm_!'1�?#            �H@        ������������������������       �                     2@        L       Q                    @D@��� ��?             ?@        M       P                   `n@�q�q�?             @        N       O                    a@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        R       W                   �d@HP�s��?             9@        S       V                    @J@����X�?             @       T       U                    �H@      �?             @        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     2@        Y       Z                    �?      �?              @        ������������������������       �                      @        [       \                   `e@�q�q�?             @       ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     &@        ������������������������       �                     5@        `       �                    �?�E����?Y             b@       a       p                   pa@��]�T��?H            �^@       b       c                    �H@��a�n`�?%             O@       ������������������������       �                     ?@        d       i                   @^@�n`���?             ?@        e       f                    ]@և���X�?             @        ������������������������       �                     �?        g       h                     J@      �?             @        ������������������������       �                     @        ������������������������       �                     @        j       o                 ����?      �?             8@        k       n                    �J@���Q��?             @       l       m                    �?�q�q�?             @       ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     3@        q       v                   0d@�-ῃ�?#            �N@        r       u                    @      �?              @        s       t                   �Z@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        w       �                   �c@�#ʆA��?            �J@       x       �                    r@և���X�?            �A@       y       �                    �H@      �?             @@       z       �                    �G@�G�z��?             4@       {       |                    @C@���Q��?             .@        ������������������������       �                      @        }       �                   pb@�	j*D�?             *@       ~                           m@X�<ݚ�?             "@        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     @        �       �                   @_@�8��8��?             (@        �       �                   @c@      �?             @       �       �                   �o@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     2@        �       �                   �Y@���N8�?             5@        ������������������������       �                     �?        ������������������������       �                     4@        �       �                    _@b�S���?�            �u@        �       �                    `@H��?"�?7             U@       �       �                   �?�g�y��?'             O@        �       �                 833�?���}<S�?             7@       �       �                    п���7�?             6@        �       �                   `]@      �?              @       ������������������������       �                     @        �       �                    �N@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     ,@        ������������������������       �                     �?        ������������������������       �                    �C@        �       �                    �O@8�A�0��?             6@       �       �                   �a@      �?             2@        �       �                   �\@      �?              @        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �?z�G�z�?             $@        ������������������������       �                     �?        �       �                   Pc@�<ݚ�?             "@        ������������������������       �                     @        �       �                    �N@      �?             @       ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     @        �       �                   �o@      �?�            �p@       �       �                 ����?+�M��?Z            �`@        �       �                    �?��.��?,            �N@        ������������������������       �                     *@        �       �                   Pd@�q�q�?$             H@       �       �                    m@�E��ӭ�?             B@       �       �                    �?z�G�z�?             >@       �       �                   �c@      �?             4@       �       �                    �L@r�q��?             2@        ������������������������       �                     @        �       �                   pb@d}h���?             ,@        ������������������������       �                     �?        �       �                   �\@8�Z$���?             *@        �       �                   Pj@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                   �\@�C��2(�?	             &@        �       �                    �N@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        �       �                 hff�?ףp=
�?             $@       ������������������������       �                      @        �       �                   �i@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �       �                    @M@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     (@        �       �                    �?d1<+�C�?.            @R@       �       �                 ����?"pc�
�?"            �K@        �       �                   ph@�X�<ݺ?             2@        �       �                     M@      �?             @        ������������������������       �                     �?        �       �                    �?�q�q�?             @       �       �                   pd@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     ,@        �       �                   �c@���"͏�?            �B@       �       �                 `ff@ףp=
�?             >@       �       �                 pff�?�nkK�?             7@        �       �                   �^@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �        	             4@        �       �                     P@����X�?             @       ������������������������       �                     @        ������������������������       �                      @        �       �                   @k@؇���X�?             @        ������������������������       �                     @        �       �                   �m@�q�q�?             @       �       �                    �L@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     2@        �                          �b@R=6�z�?R            @`@       �       �                   �a@�@��3Z�??            �X@       �       �                   Xy@�w��@�?'            �O@       �       �                 ����?j�g�y�?&             O@        �       �                   Pt@���|���?             6@       �       �                     N@�<ݚ�?             2@        �       �                    �?      �?              @        ������������������������       �                     @        �       �                    `@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     $@        ������������������������       �                     @        �       �                   Pr@�(\����?             D@       ������������������������       �                     ?@        �       �                    ^@�����H�?             "@        �       �                   �Y@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        �       �                   Hs@��?^�k�?            �A@       ������������������������       �                     7@        �       �                 ����?�8��8��?	             (@        ������������������������       �                     @        �       �                    �P@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?              
                   �?     ��?             @@             	                ���@�G�z��?
             4@                               �c@ҳ�wY;�?             1@        ������������������������       �                      @                              pff�?�q�q�?             "@                               �q@؇���X�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                     @                                �d@r�q��?	             (@                               �t@ףp=
�?             $@       ������������������������       �                     @                                d@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @                                Pe@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        �t�bh�h)h,K ��h.��R�(KMKK��h^�B0  6n����?�� ���?����=�?���
���?�|���?Y�����?h/�����?&���^B�?;�;��?vb'vb'�?      �?      �?              �?      �?      �?              �?      �?              �?                      �?S֔5eM�?���)k��?�s?�s?�?���?�;�;�?�؉�؉�?      �?        UUUUUU�?UUUUUU�?;�;��?;�;��?�$I�$I�?�m۶m��?      �?      �?              �?      �?                      �?              �?�������?�������?              �?      �?        y��x���?�!�!�?��jq��?h *�3�?�Mozӛ�?d!Y�B�?�q�q�?�q�q�?      �?                      �?      �?        I�$I�$�?n۶m۶�?UUUUUU�?�������?�7��Mo�?d!Y�B�?vb'vb'�?;�;��?      �?      �?              �?      �?              �?              �?                      �?      �?      �?�k(���?(�����?�m۶m��?�$I�$I�?333333�?�������?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?                      �?              �?      �?              �?        ;�;��?�؉�؉�?�������?�������?              �?      �?      �?      �?                      �?              �?      �?        �r
^N��??4և���?�cj`��?
qV~B��?��&�l��?6�d�M6�?>�����?	�=����?�q�q�?r�q��?      �?        �$I�$I�?�m۶m��?              �?      �?        Y�Cc�?9/���?      �?        �{����?�B!��?UUUUUU�?UUUUUU�?UUUUUU�?UUUUUU�?      �?                      �?      �?        q=
ףp�?{�G�z�?�m۶m��?�$I�$I�?      �?      �?      �?                      �?      �?              �?              �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?              �?              �?        �q�q�?r�q��?jW�v%j�?KԮD�J�?�c�1Ƹ?�s�9��?              �?�c�1��?�9�s��?۶m۶m�?�$I�$I�?              �?      �?      �?      �?                      �?      �?      �?333333�?�������?UUUUUU�?UUUUUU�?              �?      �?              �?                      �?�).�u�?�����?      �?      �?      �?      �?      �?                      �?              �?e�Cj���?5�x+��?�$I�$I�?۶m۶m�?      �?      �?�������?�������?333333�?�������?              �?vb'vb'�?;�;��?r�q��?�q�q�?              �?      �?              �?                      �?UUUUUU�?UUUUUU�?      �?      �?      �?      �?              �?      �?              �?              �?                      �?      �?        �a�a�?��y��y�?      �?                      �?��C��:�?2)^ ���?1�0��?�<��<��?�B!��?��{���?d!Y�B�?ӛ���7�?F]t�E�?�.�袋�?      �?      �?              �?      �?      �?              �?      �?                      �?      �?                      �?/�袋.�?颋.���?      �?      �?      �?      �?              �?      �?        �������?�������?              �?�q�q�?9��8���?              �?      �?      �?              �?      �?                      �?      �?      �?�n�Wc"�?�HT�n�?�����?������?      �?        UUUUUU�?�������?�q�q�?r�q��?�������?�������?      �?      �?�������?UUUUUU�?      �?        I�$I�$�?۶m۶m�?              �?;�;��?;�;��?      �?      �?              �?      �?        ]t�E�?F]t�E�?      �?      �?      �?                      �?      �?                      �?�������?�������?      �?              �?      �?              �?      �?        UUUUUU�?UUUUUU�?      �?                      �?      �?        �1bĈ�?ݹs�Ν�?F]t�E�?/�袋.�?�q�q�?��8��8�?      �?      �?              �?UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?              �?*�Y7�"�?v�)�Y7�?�������?�������?d!Y�B�?�Mozӛ�?UUUUUU�?UUUUUU�?              �?      �?                      �?�$I�$I�?�m۶m��?              �?      �?        ۶m۶m�?�$I�$I�?      �?        UUUUUU�?UUUUUU�?      �?      �?      �?                      �?      �?                      �?S+�R+��?Wj�Vj��?����>4�?���S�r�?AA�?�}��}��?��{���?B!�B�?]t�E]�?F]t�E�?9��8���?�q�q�?      �?      �?              �?�������?�������?              �?      �?              �?                      �?�������?333333�?              �?�q�q�?�q�q�?      �?      �?              �?      �?                      �?      �?        �A�A�?_�_��?              �?UUUUUU�?UUUUUU�?              �?UUUUUU�?�������?              �?      �?              �?      �?�������?�������?�������?�������?      �?        UUUUUU�?UUUUUU�?�$I�$I�?۶m۶m�?      �?                      �?      �?                      �?�������?UUUUUU�?�������?�������?      �?        UUUUUU�?UUUUUU�?              �?      �?              �?      �?              �?      �?        �t�bubhhubh)��}�(hhhhhNhKhKhG        hh%hNhJ�BHzhG        hNhG        hNhBKhDKhEh)h,K ��h.��R�(KK��h^�C              �?�t�bhQhchLC       ���R�hgKhhhkKh)h,K ��h.��R�(KK��hL�C       �t�bK��R�}�(hKhuMhvh)h,K ��h.��R�(KM��h}�B@F         �                 ����?�[��N�?�           ��@                                   I@��)��?�            �v@                                  �Z@�iʫ{�?"            �J@        ������������������������       �                     ,@                                   �?�θ�?            �C@                                  `R@      �?             8@                                  Z@����X�?             5@        ������������������������       �                      @        	       
                 ��������y4F�?             3@        ������������������������       �                      @                                    M@�t����?             1@                                hff�?�q�q�?             @                                  @F@      �?             @        ������������������������       �                     �?                                   ]@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        ������������������������       �                     &@        ������������������������       �                     @        ������������������������       �                     .@               y                   pq@�8a�ME�?�            �s@              4                   `_@�����=�?�            0p@                                  @V@�`���?            �H@        ������������������������       �                     @               )                    @L@~�4_�g�?             F@                                 �]@�n_Y�K�?             :@                                  �Y@r�q��?             @        ������������������������       �                     �?        ������������������������       �                     @                                   �X@      �?             4@        ������������������������       �                      @        !       $                   �e@r�q��?             2@        "       #                   @]@      �?             @        ������������������������       �                      @        ������������������������       �                      @        %       (                   �Y@@4և���?	             ,@        &       '                    �?�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     &@        *       3                   Xp@r�q��?             2@       +       2                    k@�t����?             1@        ,       1                   �j@�q�q�?             @       -       0                    �?z�G�z�?             @        .       /                    @N@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     &@        ������������������������       �                     �?        5       x                    �?�̐d��?w            @j@       6       w                   �e@N���X�?c            �e@       7       X                    c@Ԫ2��?b            `e@        8       =                   �\@"�W1��?.            �T@        9       <                   �m@     ��?             0@       :       ;                   �b@      �?             (@       ������������������������       �                     "@        ������������������������       �                     @        ������������������������       �                     @        >       C                    �J@6YE�t�?&            �P@       ?       @                   �a@г�wY;�?             A@       ������������������������       �                     @@        A       B                   pb@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        D       I                    �L@     ��?             @@        E       H                 ����?X�<ݚ�?             "@       F       G                   @k@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     @        J       K                    `@�㙢�c�?             7@        ������������������������       �                     @        L       U                   �o@������?
             1@       M       N                   p`@؇���X�?             ,@        ������������������������       �                     @        O       T                 ����?"pc�
�?             &@       P       Q                    �?ףp=
�?             $@       ������������������������       �                     @        R       S                   `a@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     �?        V       W                    @P@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        Y       p                 hff�?������?4            @V@       Z       ]                   �c@86��Z�?-            �S@        [       \                    b@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ^       m                    �?Х-��ٹ?*            �R@       _       f                   �[@���(-�?(            @R@        `       a                   �c@�r����?	             .@        ������������������������       �                     �?        b       e                    �?@4և���?             ,@        c       d                   �e@r�q��?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        g       l                   `@ _�@�Y�?             M@        h       i                   �o@P���Q�?             4@       ������������������������       �        
             0@        j       k                   0p@      �?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     C@        n       o                   po@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        q       v                     K@z�G�z�?             $@       r       u                   �`@�q�q�?             @       s       t                   e@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                      @        ������������������������       �                    �B@        z       �                   ``@ؓ��M{�?$            �K@       {       �                   hr@��}*_��?             ;@        |                          �q@�8��8��?             (@       }       ~                   �q@      �?             @       ������������������������       �                     @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    �?���Q��?             .@       �       �                    �L@�	j*D�?             *@       �       �                   �]@      �?              @        �       �                   (@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     @        �       �                    �M@���Q��?             @        ������������������������       �                      @        �       �                   xt@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                      @        �       �                 ����?      �?             <@       �       �                   �b@�q�q�?             8@        �       �                   Xr@�q�q�?             @        ������������������������       �                     �?        �       �                    �?z�G�z�?             @        ������������������������       �                      @        �       �                   �r@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   @g@r�q��?             2@       �       �                   �c@      �?
             0@        �       �                   �c@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     *@        ������������������������       �                      @        ������������������������       �                     @        �                         8s@ByL5���?�            �v@       �       �                   �b@PN��T'�?�            @t@       �       �                    �R@��P��i�?�            �q@       �       �                    _@	��B�?�            Pq@       �       �                 `ff@@+K&:~�?\             c@       �       �                    �Q@��ɉ�?O            @`@       �       �                    �?��v��?K            @_@       ������������������������       �        /            �R@        �       �                    �?�IєX�?            �I@       �       �                 ����?H%u��?             9@        �       �                    �L@�q�q�?             @        ������������������������       �                     �?        �       �                   �]@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                    `@�}�+r��?
             3@        ������������������������       �                     �?        ������������������������       �        	             2@        ������������������������       �                     :@        �       �                   c@z�G�z�?             @       ������������������������       �                     @        ������������������������       �                     �?        �       �                   �k@��2(&�?             6@        ������������������������       �                     $@        �       �                    @      �?             (@        ������������������������       �                     �?        �       �                   �`@"pc�
�?             &@        �       �                    �?�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                      @        �       �                   �b@Tb.��?O            @_@       �       �                    �?�_�s���?B            @Y@       �       �                    �Q@����?�?2            @T@       �       �                   P`@R���Q�?1             T@       �       �                   `@ \� ���?            �H@        �       �                    �?      �?              @        ������������������������       �                     �?        �       �                    �I@����X�?             @        ������������������������       �                      @        ������������������������       �                     @        �       �                 ���@�p ��?            �D@       �       �                 ����?�<ݚ�?             ;@       �       �                    g@؇���X�?             5@        ������������������������       �                     �?        �       �                    �?ףp=
�?             4@       �       �                 ����?�IєX�?
             1@        �       �                     G@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        ������������������������       �                     ,@        �       �                   �l@�q�q�?             @        ������������������������       �                      @        ������������������������       �                     �?        �       �                   p`@      �?             @        ������������������������       �                      @        �       �                    @J@      �?             @        ������������������������       �                      @        �       �                   a@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                     ,@        ������������������������       �                     ?@        ������������������������       �                     �?        ������������������������       �                     4@        �       �                    �?�q�q�?             8@       �       �                   pa@z�G�z�?             4@        �       �                   `c@      �?              @       �       �                    @M@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     @        ������������������������       �                     (@        ������������������������       �                     @        �       �                   `c@      �?             @        ������������������������       �                      @        ������������������������       �                      @        �       �                   �\@�K��&�?"            �E@        ������������������������       �                     @        �       �                 `ff@�G�z��?             D@       �       �                   @c@     ��?             @@        ������������������������       �                     @        �       �                 ����?l��[B��?             =@        �       �                    �K@r�q��?             @        ������������������������       �                     @        �       �                    @M@�q�q�?             @        ������������������������       �                     �?        ������������������������       �                      @        �       �                    p@\X��t�?             7@       �       �                   @j@�E��ӭ�?             2@        �       �                   �c@X�<ݚ�?             "@        ������������������������       �                     @        �       �                   �`@z�G�z�?             @        ������������������������       �                     �?        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                     @                                  @O@      �?              @       ������������������������       �                     @        ������������������������       �                     �?                                �d@�&!��?            �E@                               Ps@��%��?            �B@                                �a@����X�?             @        ������������������������       �                      @        ������������������������       �                     @                              033�?���Q��?             >@       	                        �b@
;&����?             7@       
                         T@d}h���?             ,@        ������������������������       �                     �?                                 @K@8�Z$���?             *@                                �?����X�?             @                               �Y@���Q��?             @        ������������������������       �                      @                                `]@�q�q�?             @        ������������������������       �                     �?                                  H@      �?              @        ������������������������       �                     �?        ������������������������       �                     �?        ������������������������       �                      @        ������������������������       �                     @        ������������������������       �                     "@        ������������������������       �                     @        ������������������������       �                     @        �t�bh�h)h,K ��h.��R�(KMKK��h^�B�  B~�9�J�?�@c�Z�?Np	���?d����?�琚`��?
�[���?              �?�؉�؉�?ى�؉��?      �?      �?�$I�$I�?�m۶m��?      �?        (������?6��P^C�?      �?        �?<<<<<<�?UUUUUU�?UUUUUU�?      �?      �?              �?UUUUUU�?UUUUUU�?              �?      �?                      �?              �?      �?                      �?,��O[�?�O[h���?.�!J��?F�y�b4�?և���X�?����S�?      �?        ��.���?/�袋.�?;�;��?ى�؉��?UUUUUU�?�������?      �?                      �?      �?      �?              �?�������?UUUUUU�?      �?      �?      �?                      �?n۶m۶�?�$I�$I�?UUUUUU�?UUUUUU�?      �?                      �?      �?        UUUUUU�?�������?�?<<<<<<�?UUUUUU�?UUUUUU�?�������?�������?UUUUUU�?UUUUUU�?              �?      �?                      �?      �?                      �?      �?        ��	��	�? �����?�O2�0�?_�6��<�?$���>��?p�}��?^�ڕ�]�?�ڕ�]��?      �?      �?      �?      �?      �?                      �?              �?'�l��&�?e�M6�d�?�?�?      �?              �?      �?              �?      �?              �?      �?�q�q�?r�q��?UUUUUU�?UUUUUU�?              �?      �?                      �?�7��Mo�?d!Y�B�?      �?        xxxxxx�?�?۶m۶m�?�$I�$I�?      �?        /�袋.�?F]t�E�?�������?�������?      �?        UUUUUU�?UUUUUU�?      �?                      �?              �?UUUUUU�?UUUUUU�?              �?      �?        ؽ�u�{�?B�P�"�?�Z܄��?h *�3�?      �?      �?      �?                      �?K~��K�?O贁N�?��իW��?�P�B�
�?�������?�?              �?n۶m۶�?�$I�$I�?�������?UUUUUU�?      �?                      �?      �?        #,�4�r�?�{a���?ffffff�?�������?      �?              �?      �?              �?      �?              �?              �?      �?              �?      �?        �������?�������?UUUUUU�?UUUUUU�?�������?�������?              �?      �?                      �?      �?                      �?      �?        	� O	�?�־a��?B{	�%��?_B{	�%�?UUUUUU�?UUUUUU�?      �?      �?              �?      �?                      �?333333�?�������?vb'vb'�?;�;��?      �?      �?      �?      �?      �?                      �?      �?        �������?333333�?              �?UUUUUU�?UUUUUU�?      �?                      �?              �?      �?      �?�������?�������?UUUUUU�?UUUUUU�?      �?        �������?�������?              �?UUUUUU�?UUUUUU�?              �?      �?        �������?UUUUUU�?      �?      �?UUUUUU�?UUUUUU�?      �?                      �?      �?                      �?      �?        �7PØ��?�+�U�?h/�����?&���^B�?i��ٹT�?Sm��h��?���ޓ�?�(����?Cy�5��?l(�����? �����??�?��?�~j�t��?�Zd;�?              �?�?�?���Q��?)\���(�?UUUUUU�?UUUUUU�?      �?        �������?�������?              �?      �?        (�����?�5��P�?      �?                      �?              �?�������?�������?              �?      �?        t�E]t�?��.���?              �?      �?      �?      �?        F]t�E�?/�袋.�?UUUUUU�?UUUUUU�?              �?      �?                      �?/�$��?9��v���?Q`ҩy�?��g����?�n���?~X�<��?333333�?333333�?և���X�?
^N��)�?      �?      �?      �?        �m۶m��?�$I�$I�?              �?      �?        ��+Q��?Q��+Q�?�q�q�?9��8���?�$I�$I�?۶m۶m�?      �?        �������?�������?�?�?UUUUUU�?UUUUUU�?              �?      �?                      �?UUUUUU�?UUUUUU�?              �?      �?              �?      �?              �?      �?      �?      �?              �?      �?      �?                      �?              �?              �?      �?                      �?UUUUUU�?UUUUUU�?�������?�������?      �?      �?�������?�������?              �?      �?                      �?              �?      �?              �?      �?              �?      �?        ���)k��?��)kʚ�?              �?�������?�������?      �?      �?      �?        GX�i���?���=��?UUUUUU�?�������?              �?UUUUUU�?UUUUUU�?      �?                      �?!Y�B�?��Moz��?�q�q�?r�q��?�q�q�?r�q��?              �?�������?�������?              �?      �?              �?                      �?      �?      �?              �?      �?        S֔5eM�?֔5eMY�?}���g�?���L�?�m۶m��?�$I�$I�?              �?      �?        �������?333333�?Y�B��?�Mozӛ�?۶m۶m�?I�$I�$�?      �?        ;�;��?;�;��?�$I�$I�?�m۶m��?�������?333333�?              �?UUUUUU�?UUUUUU�?      �?              �?      �?              �?      �?                      �?              �?      �?                      �?              �?�t�bubhhubehhub.